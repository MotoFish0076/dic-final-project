.SUBCKT CIM_adder_tree VSS VDD  rst_n clk Input_1[3] Input_1[2] Input_1[1] Input_1[0] Input_2[3] Input_2[2] Input_2[1] Input_2[0] Input_3[3] Input_3[2] Input_3[1] Input_3[0] Input_4[3] Input_4[2] Input_4[1] Input_4[0] Input_5[3] Input_5[2] Input_5[1] Input_5[0] Input_6[3] Input_6[2] Input_6[1] Input_6[0] Input_7[3] Input_7[2] Input_7[1] Input_7[0] Input_8[3] Input_8[2] Input_8[1] Input_8[0] Input_9[3] Input_9[2] Input_9[1] Input_9[0] Input_10[3] Input_10[2] Input_10[1] Input_10[0] Input_11[3] Input_11[2] Input_11[1] Input_11[0] Input_12[3] Input_12[2] Input_12[1] Input_12[0] Input_13[3] Input_13[2] Input_13[1] Input_13[0] Input_14[3] Input_14[2] Input_14[1] Input_14[0] Input_15[3] Input_15[2] Input_15[1] Input_15[0] Input_16[3] Input_16[2] Input_16[1] Input_16[0] Input_17[3] Input_17[2] Input_17[1] Input_17[0] Input_18[3] Input_18[2] Input_18[1] Input_18[0] Input_19[3] Input_19[2] Input_19[1] Input_19[0] Input_20[3] Input_20[2] Input_20[1] Input_20[0] Input_21[3] Input_21[2] Input_21[1] Input_21[0] Input_22[3] Input_22[2] Input_22[1] Input_22[0] Input_23[3] Input_23[2] Input_23[1] Input_23[0] Input_24[3] Input_24[2] Input_24[1] Input_24[0] Input_25[3] Input_25[2] Input_25[1] Input_25[0] Input_26[3] Input_26[2] Input_26[1] Input_26[0] Input_27[3] Input_27[2] Input_27[1] Input_27[0] Input_28[3] Input_28[2] Input_28[1] Input_28[0] Input_29[3] Input_29[2] Input_29[1] Input_29[0] Input_30[3] Input_30[2] Input_30[1] Input_30[0] Input_31[3] Input_31[2] Input_31[1] Input_31[0] Input_32[3] Input_32[2] Input_32[1] Input_32[0] out_valid Output[12] Output[11] Output[10] Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0]
XU82 VSS VDD  cnt[1] cnt[0] n149 NAND2xp5_ASAP7_75t_R
XU85 VSS VDD  cnt[2] n565 n152 NAND2xp5_ASAP7_75t_R
Xadd_123 VSS VDD  Output[12] Output[11] Output[10] Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0] n233 shift_buffer[11] shift_buffer[10] shift_buffer[9] shift_buffer[8] shift_buffer[7] shift_buffer[6] shift_buffer[5] shift_buffer[4] shift_buffer[3] shift_buffer[2] shift_buffer[1] shift_buffer[0] n233 N309 N308 N307 N306 N305 N304 N303 N302 N301 N300 N299 N298 N297 CIM_adder_tree_DW01_add_0
Xadd_0_root_add_0_root_add_96_31 VSS VDD  n233 N224 N223 N222 N221 N220 N219 N218 n167 n233 N260 N259 N258 N257 N256 N255 N254 n182 n233 N279 N278 N277 N276 N275 N274 N273 N272 N271 CIM_adder_tree_DW01_add_1
Xadd_1_root_add_0_root_add_96_31_U1_1 VSS VDD  add_1_root_add_0_root_add_96_31_A_1_ add_1_root_add_0_root_add_96_31_B_1_ n165 n533 n532 FAx1_ASAP7_75t_R
Xadd_1_root_add_0_root_add_96_31_U1_2 VSS VDD  add_1_root_add_0_root_add_96_31_A_2_ add_1_root_add_0_root_add_96_31_B_2_ n544 n535 n534 FAx1_ASAP7_75t_R
Xadd_1_root_add_0_root_add_96_31_U1_3 VSS VDD  add_1_root_add_0_root_add_96_31_A_3_ add_1_root_add_0_root_add_96_31_B_3_ n545 n537 n536 FAx1_ASAP7_75t_R
Xadd_1_root_add_0_root_add_96_31_U1_4 VSS VDD  add_1_root_add_0_root_add_96_31_A_4_ add_1_root_add_0_root_add_96_31_B_4_ n546 n539 n538 FAx1_ASAP7_75t_R
Xadd_1_root_add_0_root_add_96_31_U1_5 VSS VDD  add_1_root_add_0_root_add_96_31_A_5_ add_1_root_add_0_root_add_96_31_B_5_ n547 n541 n540 FAx1_ASAP7_75t_R
Xadd_1_root_add_0_root_add_96_31_U1_6 VSS VDD  add_1_root_add_0_root_add_96_31_A_6_ add_1_root_add_0_root_add_96_31_B_6_ n548 n543 n542 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_1 VSS VDD  N155 N146 n166 n516 n515 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_2 VSS VDD  N156 N147 n527 n518 n517 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_3 VSS VDD  N157 N148 n528 n520 n519 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_4 VSS VDD  N158 N149 n529 n522 n521 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_5 VSS VDD  N159 N150 n530 n524 n523 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_6 VSS VDD  N160 N151 n531 n526 n525 FAx1_ASAP7_75t_R
Xadd_6_root_add_0_root_add_96_31_U1_1 VSS VDD  N47 add_6_root_add_0_root_add_96_31_B_1_ n164 n502 n501 FAx1_ASAP7_75t_R
Xadd_6_root_add_0_root_add_96_31_U1_2 VSS VDD  N48 add_6_root_add_0_root_add_96_31_B_2_ n511 n504 n503 FAx1_ASAP7_75t_R
Xadd_6_root_add_0_root_add_96_31_U1_3 VSS VDD  N49 add_6_root_add_0_root_add_96_31_B_3_ n512 n506 n505 FAx1_ASAP7_75t_R
Xadd_6_root_add_0_root_add_96_31_U1_4 VSS VDD  N50 add_6_root_add_0_root_add_96_31_B_4_ n513 n508 n507 FAx1_ASAP7_75t_R
Xadd_6_root_add_0_root_add_96_31_U1_5 VSS VDD  N51 add_6_root_add_0_root_add_96_31_B_5_ n514 n510 n509 FAx1_ASAP7_75t_R
Xadd_3_root_add_0_root_add_96_31_U1_1 VSS VDD  N56 N38 n163 n488 n487 FAx1_ASAP7_75t_R
Xadd_3_root_add_0_root_add_96_31_U1_2 VSS VDD  N57 N39 n497 n490 n489 FAx1_ASAP7_75t_R
Xadd_3_root_add_0_root_add_96_31_U1_3 VSS VDD  N58 N40 n498 n492 n491 FAx1_ASAP7_75t_R
Xadd_3_root_add_0_root_add_96_31_U1_4 VSS VDD  N59 N41 n499 n494 n493 FAx1_ASAP7_75t_R
Xadd_3_root_add_0_root_add_96_31_U1_5 VSS VDD  N60 N42 n500 n496 n495 FAx1_ASAP7_75t_R
Xadd_14_root_add_0_root_add_96_31_U1_1 VSS VDD  N128 N65 n158 n477 n476 FAx1_ASAP7_75t_R
Xadd_14_root_add_0_root_add_96_31_U1_2 VSS VDD  N129 N66 n484 n479 n478 FAx1_ASAP7_75t_R
Xadd_14_root_add_0_root_add_96_31_U1_3 VSS VDD  N130 N67 n485 n481 n480 FAx1_ASAP7_75t_R
Xadd_14_root_add_0_root_add_96_31_U1_4 VSS VDD  N131 N68 n486 n483 n482 FAx1_ASAP7_75t_R
Xadd_15_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_15[1] Input_14[1] n197 n469 n468 FAx1_ASAP7_75t_R
Xadd_15_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_15[2] Input_14[2] n474 n471 n470 FAx1_ASAP7_75t_R
Xadd_15_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_15[3] Input_14[3] n475 n473 n472 FAx1_ASAP7_75t_R
Xadd_29_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_30[1] Input_2[1] n193 n461 n460 FAx1_ASAP7_75t_R
Xadd_29_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_30[2] Input_2[2] n466 n463 n462 FAx1_ASAP7_75t_R
Xadd_29_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_30[3] Input_2[3] n467 n465 n464 FAx1_ASAP7_75t_R
Xadd_12_root_add_0_root_add_96_31_U1_1 VSS VDD  N200 N236 n157 n450 n449 FAx1_ASAP7_75t_R
Xadd_12_root_add_0_root_add_96_31_U1_2 VSS VDD  N201 N237 n457 n452 n451 FAx1_ASAP7_75t_R
Xadd_12_root_add_0_root_add_96_31_U1_3 VSS VDD  N202 N238 n458 n454 n453 FAx1_ASAP7_75t_R
Xadd_12_root_add_0_root_add_96_31_U1_4 VSS VDD  N203 N239 n459 n456 n455 FAx1_ASAP7_75t_R
Xadd_17_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_12[1] Input_6[1] n196 n442 n441 FAx1_ASAP7_75t_R
Xadd_17_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_12[2] Input_6[2] n447 n444 n443 FAx1_ASAP7_75t_R
Xadd_17_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_12[3] Input_6[3] n448 n446 n445 FAx1_ASAP7_75t_R
Xadd_25_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_26[1] Input_17[1] n192 n434 n433 FAx1_ASAP7_75t_R
Xadd_25_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_26[2] Input_17[2] n439 n436 n435 FAx1_ASAP7_75t_R
Xadd_25_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_26[3] Input_17[3] n440 n438 n437 FAx1_ASAP7_75t_R
Xadd_11_root_add_0_root_add_96_31_U1_1 VSS VDD  N110 N182 n160 n423 n422 FAx1_ASAP7_75t_R
Xadd_11_root_add_0_root_add_96_31_U1_2 VSS VDD  N111 N183 n430 n425 n424 FAx1_ASAP7_75t_R
Xadd_11_root_add_0_root_add_96_31_U1_3 VSS VDD  N112 N184 n431 n427 n426 FAx1_ASAP7_75t_R
Xadd_11_root_add_0_root_add_96_31_U1_4 VSS VDD  N113 N185 n432 n429 n428 FAx1_ASAP7_75t_R
Xadd_18_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_3[1] Input_21[1] n199 n415 n414 FAx1_ASAP7_75t_R
Xadd_18_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_3[2] Input_21[2] n420 n417 n416 FAx1_ASAP7_75t_R
Xadd_18_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_3[3] Input_21[3] n421 n419 n418 FAx1_ASAP7_75t_R
Xadd_26_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_27[1] Input_16[1] n195 n407 n406 FAx1_ASAP7_75t_R
Xadd_26_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_27[2] Input_16[2] n412 n409 n408 FAx1_ASAP7_75t_R
Xadd_26_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_27[3] Input_16[3] n413 n411 n410 FAx1_ASAP7_75t_R
Xadd_7_root_add_0_root_add_96_31_U1_1 VSS VDD  N209 N119 n159 n396 n395 FAx1_ASAP7_75t_R
Xadd_7_root_add_0_root_add_96_31_U1_2 VSS VDD  N210 N120 n403 n398 n397 FAx1_ASAP7_75t_R
Xadd_7_root_add_0_root_add_96_31_U1_3 VSS VDD  N211 N121 n404 n400 n399 FAx1_ASAP7_75t_R
Xadd_7_root_add_0_root_add_96_31_U1_4 VSS VDD  N212 N122 n405 n402 n401 FAx1_ASAP7_75t_R
Xadd_27_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_28[1] Input_8[1] n198 n388 n387 FAx1_ASAP7_75t_R
Xadd_27_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_28[2] Input_8[2] n393 n390 n389 FAx1_ASAP7_75t_R
Xadd_27_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_28[3] Input_8[3] n394 n392 n391 FAx1_ASAP7_75t_R
Xadd_28_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_29[1] Input_4[1] n194 n380 n379 FAx1_ASAP7_75t_R
Xadd_28_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_29[2] Input_4[2] n385 n382 n381 FAx1_ASAP7_75t_R
Xadd_28_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_29[3] Input_4[3] n386 n384 n383 FAx1_ASAP7_75t_R
Xadd_5_root_add_0_root_add_96_31_U1_1 VSS VDD  N173 add_5_root_add_0_root_add_96_31_B_1_ n161 n366 n365 FAx1_ASAP7_75t_R
Xadd_5_root_add_0_root_add_96_31_U1_2 VSS VDD  N174 add_5_root_add_0_root_add_96_31_B_2_ n375 n368 n367 FAx1_ASAP7_75t_R
Xadd_5_root_add_0_root_add_96_31_U1_3 VSS VDD  N175 add_5_root_add_0_root_add_96_31_B_3_ n376 n370 n369 FAx1_ASAP7_75t_R
Xadd_5_root_add_0_root_add_96_31_U1_4 VSS VDD  N176 add_5_root_add_0_root_add_96_31_B_4_ n377 n372 n371 FAx1_ASAP7_75t_R
Xadd_5_root_add_0_root_add_96_31_U1_5 VSS VDD  N177 add_5_root_add_0_root_add_96_31_B_5_ n378 n374 n373 FAx1_ASAP7_75t_R
Xadd_8_root_add_0_root_add_96_31_U1_1 VSS VDD  N137 N74 n156 n355 n354 FAx1_ASAP7_75t_R
Xadd_8_root_add_0_root_add_96_31_U1_2 VSS VDD  N138 N75 n362 n357 n356 FAx1_ASAP7_75t_R
Xadd_8_root_add_0_root_add_96_31_U1_3 VSS VDD  N139 N76 n363 n359 n358 FAx1_ASAP7_75t_R
Xadd_8_root_add_0_root_add_96_31_U1_4 VSS VDD  N140 N77 n364 n361 n360 FAx1_ASAP7_75t_R
Xadd_19_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_31[1] Input_11[1] n191 n347 n346 FAx1_ASAP7_75t_R
Xadd_19_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_31[2] Input_11[2] n352 n349 n348 FAx1_ASAP7_75t_R
Xadd_19_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_31[3] Input_11[3] n353 n351 n350 FAx1_ASAP7_75t_R
Xadd_30_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_1[1] Input_32[1] n187 n339 n338 FAx1_ASAP7_75t_R
Xadd_30_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_1[2] Input_32[2] n344 n341 n340 FAx1_ASAP7_75t_R
Xadd_30_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_1[3] Input_32[3] n345 n343 n342 FAx1_ASAP7_75t_R
Xadd_13_root_add_0_root_add_96_31_U1_1 VSS VDD  N245 N263 n154 n328 n327 FAx1_ASAP7_75t_R
Xadd_13_root_add_0_root_add_96_31_U1_2 VSS VDD  N246 N264 n335 n330 n329 FAx1_ASAP7_75t_R
Xadd_13_root_add_0_root_add_96_31_U1_3 VSS VDD  N247 N265 n336 n332 n331 FAx1_ASAP7_75t_R
Xadd_13_root_add_0_root_add_96_31_U1_4 VSS VDD  N248 N266 n337 n334 n333 FAx1_ASAP7_75t_R
Xadd_16_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_7[1] Input_13[1] n189 n320 n319 FAx1_ASAP7_75t_R
Xadd_16_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_7[2] Input_13[2] n325 n322 n321 FAx1_ASAP7_75t_R
Xadd_16_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_7[3] Input_13[3] n326 n324 n323 FAx1_ASAP7_75t_R
Xadd_24_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_25[1] Input_9[1] n185 n312 n311 FAx1_ASAP7_75t_R
Xadd_24_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_25[2] Input_9[2] n317 n314 n313 FAx1_ASAP7_75t_R
Xadd_24_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_25[3] Input_9[3] n318 n316 n315 FAx1_ASAP7_75t_R
Xadd_4_root_add_0_root_add_96_31_U1_1 VSS VDD  N164 N227 n162 n298 n297 FAx1_ASAP7_75t_R
Xadd_4_root_add_0_root_add_96_31_U1_2 VSS VDD  N165 N228 n307 n300 n299 FAx1_ASAP7_75t_R
Xadd_4_root_add_0_root_add_96_31_U1_3 VSS VDD  N166 N229 n308 n302 n301 FAx1_ASAP7_75t_R
Xadd_4_root_add_0_root_add_96_31_U1_4 VSS VDD  N167 N230 n309 n304 n303 FAx1_ASAP7_75t_R
Xadd_4_root_add_0_root_add_96_31_U1_5 VSS VDD  N168 N231 n310 n306 n305 FAx1_ASAP7_75t_R
Xadd_9_root_add_0_root_add_96_31_U1_1 VSS VDD  N83 N101 n155 n287 n286 FAx1_ASAP7_75t_R
Xadd_9_root_add_0_root_add_96_31_U1_2 VSS VDD  N84 N102 n294 n289 n288 FAx1_ASAP7_75t_R
Xadd_9_root_add_0_root_add_96_31_U1_3 VSS VDD  N85 N103 n295 n291 n290 FAx1_ASAP7_75t_R
Xadd_9_root_add_0_root_add_96_31_U1_4 VSS VDD  N86 N104 n296 n293 n292 FAx1_ASAP7_75t_R
Xadd_23_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_24[1] Input_18[1] n190 n279 n278 FAx1_ASAP7_75t_R
Xadd_23_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_24[2] Input_18[2] n284 n281 n280 FAx1_ASAP7_75t_R
Xadd_23_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_24[3] Input_18[3] n285 n283 n282 FAx1_ASAP7_75t_R
Xadd_20_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_10[1] Input_20[1] n186 n271 n270 FAx1_ASAP7_75t_R
Xadd_20_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_10[2] Input_20[2] n276 n273 n272 FAx1_ASAP7_75t_R
Xadd_20_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_10[3] Input_20[3] n277 n275 n274 FAx1_ASAP7_75t_R
Xadd_10_root_add_0_root_add_96_31_U1_1 VSS VDD  N92 N191 n153 n260 n259 FAx1_ASAP7_75t_R
Xadd_10_root_add_0_root_add_96_31_U1_2 VSS VDD  N93 N192 n267 n262 n261 FAx1_ASAP7_75t_R
Xadd_10_root_add_0_root_add_96_31_U1_3 VSS VDD  N94 N193 n268 n264 n263 FAx1_ASAP7_75t_R
Xadd_10_root_add_0_root_add_96_31_U1_4 VSS VDD  N95 N194 n269 n266 n265 FAx1_ASAP7_75t_R
Xadd_21_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_22[1] Input_5[1] n188 n252 n251 FAx1_ASAP7_75t_R
Xadd_21_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_22[2] Input_5[2] n257 n254 n253 FAx1_ASAP7_75t_R
Xadd_21_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_22[3] Input_5[3] n258 n256 n255 FAx1_ASAP7_75t_R
Xadd_22_root_add_0_root_add_96_31_U1_1 VSS VDD  Input_23[1] Input_19[1] n184 n244 n243 FAx1_ASAP7_75t_R
Xadd_22_root_add_0_root_add_96_31_U1_2 VSS VDD  Input_23[2] Input_19[2] n249 n246 n245 FAx1_ASAP7_75t_R
Xadd_22_root_add_0_root_add_96_31_U1_3 VSS VDD  Input_23[3] Input_19[3] n250 n248 n247 FAx1_ASAP7_75t_R
Xcnt_reg_0_ VSS VDD  n240 clk n233 n558 cnt[0] ASYNC_DFFHx1_ASAP7_75t_R
Xcnt_reg_2_ VSS VDD  n563 clk n233 n558 cnt[2] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_2_ VSS VDD  n232 clk n558 n233 Output[2] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_1_ VSS VDD  n231 clk n558 n233 Output[1] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_0_ VSS VDD  n183 clk n558 n233 Output[0] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_3_ VSS VDD  n230 clk n558 n233 Output[3] ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg VSS VDD  n564 clk n558 n233 out_valid ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_4_ VSS VDD  n228 clk n558 n233 Output[4] ASYNC_DFFHx1_ASAP7_75t_R
Xcnt_reg_1_ VSS VDD  n229 clk n558 n233 cnt[1] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_5_ VSS VDD  n227 clk n558 n233 Output[5] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_6_ VSS VDD  n226 clk n558 n233 Output[6] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_3_ VSS VDD  n239 clk n558 n233 shift_buffer[3] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_2_ VSS VDD  n238 clk n558 n233 shift_buffer[2] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_1_ VSS VDD  n237 clk n558 n233 shift_buffer[1] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_0_ VSS VDD  n236 clk n558 n233 shift_buffer[0] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_5_ VSS VDD  n235 clk n558 n233 shift_buffer[5] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_4_ VSS VDD  n234 clk n558 n233 shift_buffer[4] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_7_ VSS VDD  n225 clk n558 n233 Output[7] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_11_ VSS VDD  n224 clk n558 n233 shift_buffer[11] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_10_ VSS VDD  n223 clk n558 n233 shift_buffer[10] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_9_ VSS VDD  n222 clk n558 n233 shift_buffer[9] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_8_ VSS VDD  n221 clk n558 n233 shift_buffer[8] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_7_ VSS VDD  n220 clk n558 n233 shift_buffer[7] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_6_ VSS VDD  n219 clk n558 n233 shift_buffer[6] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_8_ VSS VDD  n218 clk n558 n233 Output[8] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_9_ VSS VDD  n217 clk n558 n233 Output[9] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_10_ VSS VDD  n216 clk n558 n233 Output[10] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_11_ VSS VDD  n215 clk n558 n233 Output[11] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_12_ VSS VDD  n214 clk n558 n233 Output[12] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_0_ VSS VDD  n557 clk n558 n233 input_buffer[0] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_1_ VSS VDD  n556 clk n558 n233 input_buffer[1] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_2_ VSS VDD  n555 clk n558 n233 input_buffer[2] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_3_ VSS VDD  n554 clk n558 n233 input_buffer[3] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_4_ VSS VDD  n553 clk n558 n233 input_buffer[4] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_5_ VSS VDD  n552 clk n558 n233 input_buffer[5] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_6_ VSS VDD  n551 clk n558 n233 input_buffer[6] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_8_ VSS VDD  n549 clk n558 n233 input_buffer[8] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_7_ VSS VDD  n550 clk n558 n233 input_buffer[7] ASYNC_DFFHx1_ASAP7_75t_R
XU106 VSS VDD  n233 TIELOx1_ASAP7_75t_R
XU107 VSS VDD  n242 n625 n603 NOR2xp33_ASAP7_75t_R
XU108 VSS VDD  n242 n628 n610 NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  n169 n201 n153 AND2x2_ASAP7_75t_R
XU110 VSS VDD  n168 n200 n154 AND2x2_ASAP7_75t_R
XU111 VSS VDD  n171 n203 n155 AND2x2_ASAP7_75t_R
XU112 VSS VDD  n170 n202 n156 AND2x2_ASAP7_75t_R
XU113 VSS VDD  n173 n205 n157 AND2x2_ASAP7_75t_R
XU114 VSS VDD  n172 n204 n158 AND2x2_ASAP7_75t_R
XU115 VSS VDD  n175 n207 n159 AND2x2_ASAP7_75t_R
XU116 VSS VDD  n174 n206 n160 AND2x2_ASAP7_75t_R
XU117 VSS VDD  n176 n208 n161 AND2x2_ASAP7_75t_R
XU118 VSS VDD  n177 n209 n162 AND2x2_ASAP7_75t_R
XU119 VSS VDD  n178 n210 n163 AND2x2_ASAP7_75t_R
XU120 VSS VDD  n179 n211 n164 AND2x2_ASAP7_75t_R
XU121 VSS VDD  n180 n212 n165 AND2x2_ASAP7_75t_R
XU122 VSS VDD  n181 n213 n166 AND2x2_ASAP7_75t_R
XU123 VSS VDD  n181 n213 n167 XOR2xp5_ASAP7_75t_R
XU124 VSS VDD  Input_25[0] Input_9[0] n168 XOR2xp5_ASAP7_75t_R
XU125 VSS VDD  Input_23[0] Input_19[0] n169 XOR2xp5_ASAP7_75t_R
XU126 VSS VDD  Input_1[0] Input_32[0] n170 XOR2xp5_ASAP7_75t_R
XU127 VSS VDD  Input_10[0] Input_20[0] n171 XOR2xp5_ASAP7_75t_R
XU128 VSS VDD  Input_30[0] Input_2[0] n172 XOR2xp5_ASAP7_75t_R
XU129 VSS VDD  Input_26[0] Input_17[0] n173 XOR2xp5_ASAP7_75t_R
XU130 VSS VDD  Input_27[0] Input_16[0] n174 XOR2xp5_ASAP7_75t_R
XU131 VSS VDD  Input_29[0] Input_4[0] n175 XOR2xp5_ASAP7_75t_R
XU132 VSS VDD  n168 n200 n176 XOR2xp5_ASAP7_75t_R
XU133 VSS VDD  n169 n201 n177 XOR2xp5_ASAP7_75t_R
XU134 VSS VDD  n172 n204 n178 XOR2xp5_ASAP7_75t_R
XU135 VSS VDD  n173 n205 n179 XOR2xp5_ASAP7_75t_R
XU136 VSS VDD  n177 n209 n180 XOR2xp5_ASAP7_75t_R
XU137 VSS VDD  n179 n211 n181 XOR2xp5_ASAP7_75t_R
XU138 VSS VDD  n180 n212 n182 XOR2xp5_ASAP7_75t_R
XU139 VSS VDD  N297 n150 n183 NAND2xp5_ASAP7_75t_R
XU140 VSS VDD  Input_23[0] Input_19[0] n184 AND2x2_ASAP7_75t_R
XU141 VSS VDD  Input_25[0] Input_9[0] n185 AND2x2_ASAP7_75t_R
XU142 VSS VDD  Input_10[0] Input_20[0] n186 AND2x2_ASAP7_75t_R
XU143 VSS VDD  Input_1[0] Input_32[0] n187 AND2x2_ASAP7_75t_R
XU144 VSS VDD  Input_22[0] Input_5[0] n188 AND2x2_ASAP7_75t_R
XU145 VSS VDD  Input_7[0] Input_13[0] n189 AND2x2_ASAP7_75t_R
XU146 VSS VDD  Input_24[0] Input_18[0] n190 AND2x2_ASAP7_75t_R
XU147 VSS VDD  Input_31[0] Input_11[0] n191 AND2x2_ASAP7_75t_R
XU148 VSS VDD  Input_26[0] Input_17[0] n192 AND2x2_ASAP7_75t_R
XU149 VSS VDD  Input_30[0] Input_2[0] n193 AND2x2_ASAP7_75t_R
XU150 VSS VDD  Input_29[0] Input_4[0] n194 AND2x2_ASAP7_75t_R
XU151 VSS VDD  Input_27[0] Input_16[0] n195 AND2x2_ASAP7_75t_R
XU152 VSS VDD  Input_12[0] Input_6[0] n196 AND2x2_ASAP7_75t_R
XU153 VSS VDD  Input_15[0] Input_14[0] n197 AND2x2_ASAP7_75t_R
XU154 VSS VDD  Input_28[0] Input_8[0] n198 AND2x2_ASAP7_75t_R
XU155 VSS VDD  Input_3[0] Input_21[0] n199 AND2x2_ASAP7_75t_R
XU156 VSS VDD  Input_7[0] Input_13[0] n200 XOR2xp5_ASAP7_75t_R
XU157 VSS VDD  Input_22[0] Input_5[0] n201 XOR2xp5_ASAP7_75t_R
XU158 VSS VDD  Input_31[0] Input_11[0] n202 XOR2xp5_ASAP7_75t_R
XU159 VSS VDD  Input_24[0] Input_18[0] n203 XOR2xp5_ASAP7_75t_R
XU160 VSS VDD  Input_15[0] Input_14[0] n204 XOR2xp5_ASAP7_75t_R
XU161 VSS VDD  Input_12[0] Input_6[0] n205 XOR2xp5_ASAP7_75t_R
XU162 VSS VDD  Input_3[0] Input_21[0] n206 XOR2xp5_ASAP7_75t_R
XU163 VSS VDD  Input_28[0] Input_8[0] n207 XOR2xp5_ASAP7_75t_R
XU164 VSS VDD  n170 n202 n208 XOR2xp5_ASAP7_75t_R
XU165 VSS VDD  n171 n203 n209 XOR2xp5_ASAP7_75t_R
XU166 VSS VDD  n174 n206 n210 XOR2xp5_ASAP7_75t_R
XU167 VSS VDD  n175 n207 n211 XOR2xp5_ASAP7_75t_R
XU168 VSS VDD  n176 n208 n212 XOR2xp5_ASAP7_75t_R
XU169 VSS VDD  n178 n210 n213 XOR2xp5_ASAP7_75t_R
XU170 VSS VDD  N309 n150 n214 NAND2xp5_ASAP7_75t_R
XU171 VSS VDD  N308 n150 n215 NAND2xp5_ASAP7_75t_R
XU172 VSS VDD  N307 n150 n216 NAND2xp5_ASAP7_75t_R
XU173 VSS VDD  N306 n150 n217 NAND2xp5_ASAP7_75t_R
XU174 VSS VDD  N305 n150 n218 NAND2xp5_ASAP7_75t_R
XU175 VSS VDD  n241 n615 n614 n219 OR3x1_ASAP7_75t_R
XU176 VSS VDD  n241 n619 n618 n220 OR3x1_ASAP7_75t_R
XU177 VSS VDD  n241 n627 n626 n221 OR3x1_ASAP7_75t_R
XU178 VSS VDD  n241 n635 n634 n222 OR3x1_ASAP7_75t_R
XU179 VSS VDD  n241 n576 n575 n223 OR3x1_ASAP7_75t_R
XU180 VSS VDD  n241 n585 n584 n224 OR3x1_ASAP7_75t_R
XU181 VSS VDD  N304 n150 n225 NAND2xp5_ASAP7_75t_R
XU182 VSS VDD  N303 n150 n226 NAND2xp5_ASAP7_75t_R
XU183 VSS VDD  N302 n150 n227 NAND2xp5_ASAP7_75t_R
XU184 VSS VDD  N301 n150 n228 NAND2xp5_ASAP7_75t_R
XU185 VSS VDD  n564 N6 n229 NAND2xp5_ASAP7_75t_R
XU186 VSS VDD  N300 n150 n230 NAND2xp5_ASAP7_75t_R
XU187 VSS VDD  N298 n150 n231 NAND2xp5_ASAP7_75t_R
XU188 VSS VDD  N299 n150 n232 NAND2xp5_ASAP7_75t_R
XU189 VSS VDD  n242 n612 n615 NOR2xp33_ASAP7_75t_R
XU190 VSS VDD  n613 n563 n614 NOR2xp33_ASAP7_75t_R
XU191 VSS VDD  n242 n616 n619 NOR2xp33_ASAP7_75t_R
XU192 VSS VDD  n617 n563 n618 NOR2xp33_ASAP7_75t_R
XU193 VSS VDD  n242 n624 n627 NOR2xp33_ASAP7_75t_R
XU194 VSS VDD  n625 n563 n626 NOR2xp33_ASAP7_75t_R
XU195 VSS VDD  n242 n583 n584 NOR2xp33_ASAP7_75t_R
XU196 VSS VDD  n616 n563 n585 NOR2xp33_ASAP7_75t_R
XU197 VSS VDD  n242 n633 n634 NOR2xp33_ASAP7_75t_R
XU198 VSS VDD  n628 n563 n635 NOR2xp33_ASAP7_75t_R
XU199 VSS VDD  n242 n574 n575 NOR2xp33_ASAP7_75t_R
XU200 VSS VDD  n612 n563 n576 NOR2xp33_ASAP7_75t_R
XU201 VSS VDD  n241 n604 n603 n234 OR3x1_ASAP7_75t_R
XU202 VSS VDD  n241 n611 n610 n235 OR3x1_ASAP7_75t_R
XU203 VSS VDD  n598 n241 n242 n236 OR3x1_ASAP7_75t_R
XU204 VSS VDD  n605 n241 n242 n237 OR3x1_ASAP7_75t_R
XU205 VSS VDD  n560 n241 n242 n238 OR3x1_ASAP7_75t_R
XU206 VSS VDD  n559 n241 n242 n239 OR3x1_ASAP7_75t_R
XU207 VSS VDD  N6 n562 INVx1_ASAP7_75t_R
XU208 VSS VDD  n632 n631 n633 NOR2xp33_ASAP7_75t_R
XU209 VSS VDD  n562 n630 n631 NOR2xp33_ASAP7_75t_R
XU210 VSS VDD  n623 n622 n624 NOR2xp33_ASAP7_75t_R
XU211 VSS VDD  N6 n620 n623 NOR2xp33_ASAP7_75t_R
XU212 VSS VDD  n562 n621 n622 NOR2xp33_ASAP7_75t_R
XU213 VSS VDD  n562 n629 n583 NOR2xp33_ASAP7_75t_R
XU214 VSS VDD  cnt[1] cnt[0] n151 NOR2xp33_ASAP7_75t_R
XU215 VSS VDD  N284 n241 HB1xp67_ASAP7_75t_R
XU216 VSS VDD  n565 cnt[2] N284 NOR2xp33_ASAP7_75t_R
XU217 VSS VDD  N7 n242 HB1xp67_ASAP7_75t_R
XU218 VSS VDD  n564 n152 N7 NAND2xp5_ASAP7_75t_R
XU219 VSS VDD  n565 n149 N6 NAND2xp5_ASAP7_75t_R
XU220 VSS VDD  cnt[0] n241 n240 OR2x2_ASAP7_75t_R
XU221 VSS VDD  cnt[0] n561 INVx1_ASAP7_75t_R
XU222 VSS VDD  cnt[2] n151 n150 NAND2xp5_ASAP7_75t_R
XU223 VSS VDD  n243 N92 INVx1_ASAP7_75t_R
XU224 VSS VDD  n245 N93 INVx1_ASAP7_75t_R
XU225 VSS VDD  n247 N94 INVx1_ASAP7_75t_R
XU226 VSS VDD  n248 N95 INVx1_ASAP7_75t_R
XU227 VSS VDD  n244 n249 INVx1_ASAP7_75t_R
XU228 VSS VDD  n246 n250 INVx1_ASAP7_75t_R
XU229 VSS VDD  n251 N191 INVx1_ASAP7_75t_R
XU230 VSS VDD  n253 N192 INVx1_ASAP7_75t_R
XU231 VSS VDD  n255 N193 INVx1_ASAP7_75t_R
XU232 VSS VDD  n256 N194 INVx1_ASAP7_75t_R
XU233 VSS VDD  n252 n257 INVx1_ASAP7_75t_R
XU234 VSS VDD  n254 n258 INVx1_ASAP7_75t_R
XU235 VSS VDD  n259 N164 INVx1_ASAP7_75t_R
XU236 VSS VDD  n261 N165 INVx1_ASAP7_75t_R
XU237 VSS VDD  n263 N166 INVx1_ASAP7_75t_R
XU238 VSS VDD  n265 N167 INVx1_ASAP7_75t_R
XU239 VSS VDD  n266 N168 INVx1_ASAP7_75t_R
XU240 VSS VDD  n260 n267 INVx1_ASAP7_75t_R
XU241 VSS VDD  n262 n268 INVx1_ASAP7_75t_R
XU242 VSS VDD  n264 n269 INVx1_ASAP7_75t_R
XU243 VSS VDD  n270 N83 INVx1_ASAP7_75t_R
XU244 VSS VDD  n272 N84 INVx1_ASAP7_75t_R
XU245 VSS VDD  n274 N85 INVx1_ASAP7_75t_R
XU246 VSS VDD  n275 N86 INVx1_ASAP7_75t_R
XU247 VSS VDD  n271 n276 INVx1_ASAP7_75t_R
XU248 VSS VDD  n273 n277 INVx1_ASAP7_75t_R
XU249 VSS VDD  n278 N101 INVx1_ASAP7_75t_R
XU250 VSS VDD  n280 N102 INVx1_ASAP7_75t_R
XU251 VSS VDD  n282 N103 INVx1_ASAP7_75t_R
XU252 VSS VDD  n283 N104 INVx1_ASAP7_75t_R
XU253 VSS VDD  n279 n284 INVx1_ASAP7_75t_R
XU254 VSS VDD  n281 n285 INVx1_ASAP7_75t_R
XU255 VSS VDD  n286 N227 INVx1_ASAP7_75t_R
XU256 VSS VDD  n288 N228 INVx1_ASAP7_75t_R
XU257 VSS VDD  n290 N229 INVx1_ASAP7_75t_R
XU258 VSS VDD  n292 N230 INVx1_ASAP7_75t_R
XU259 VSS VDD  n293 N231 INVx1_ASAP7_75t_R
XU260 VSS VDD  n287 n294 INVx1_ASAP7_75t_R
XU261 VSS VDD  n289 n295 INVx1_ASAP7_75t_R
XU262 VSS VDD  n291 n296 INVx1_ASAP7_75t_R
XU263 VSS VDD  n297 add_1_root_add_0_root_add_96_31_A_1_ INVx1_ASAP7_75t_R
XU264 VSS VDD  n299 add_1_root_add_0_root_add_96_31_A_2_ INVx1_ASAP7_75t_R
XU265 VSS VDD  n301 add_1_root_add_0_root_add_96_31_A_3_ INVx1_ASAP7_75t_R
XU266 VSS VDD  n303 add_1_root_add_0_root_add_96_31_A_4_ INVx1_ASAP7_75t_R
XU267 VSS VDD  n305 add_1_root_add_0_root_add_96_31_A_5_ INVx1_ASAP7_75t_R
XU268 VSS VDD  n306 add_1_root_add_0_root_add_96_31_A_6_ INVx1_ASAP7_75t_R
XU269 VSS VDD  n298 n307 INVx1_ASAP7_75t_R
XU270 VSS VDD  n300 n308 INVx1_ASAP7_75t_R
XU271 VSS VDD  n302 n309 INVx1_ASAP7_75t_R
XU272 VSS VDD  n304 n310 INVx1_ASAP7_75t_R
XU273 VSS VDD  n311 N245 INVx1_ASAP7_75t_R
XU274 VSS VDD  n313 N246 INVx1_ASAP7_75t_R
XU275 VSS VDD  n315 N247 INVx1_ASAP7_75t_R
XU276 VSS VDD  n316 N248 INVx1_ASAP7_75t_R
XU277 VSS VDD  n312 n317 INVx1_ASAP7_75t_R
XU278 VSS VDD  n314 n318 INVx1_ASAP7_75t_R
XU279 VSS VDD  n319 N263 INVx1_ASAP7_75t_R
XU280 VSS VDD  n321 N264 INVx1_ASAP7_75t_R
XU281 VSS VDD  n323 N265 INVx1_ASAP7_75t_R
XU282 VSS VDD  n324 N266 INVx1_ASAP7_75t_R
XU283 VSS VDD  n320 n325 INVx1_ASAP7_75t_R
XU284 VSS VDD  n322 n326 INVx1_ASAP7_75t_R
XU285 VSS VDD  n327 N173 INVx1_ASAP7_75t_R
XU286 VSS VDD  n329 N174 INVx1_ASAP7_75t_R
XU287 VSS VDD  n331 N175 INVx1_ASAP7_75t_R
XU288 VSS VDD  n333 N176 INVx1_ASAP7_75t_R
XU289 VSS VDD  n334 N177 INVx1_ASAP7_75t_R
XU290 VSS VDD  n328 n335 INVx1_ASAP7_75t_R
XU291 VSS VDD  n330 n336 INVx1_ASAP7_75t_R
XU292 VSS VDD  n332 n337 INVx1_ASAP7_75t_R
XU293 VSS VDD  n338 N137 INVx1_ASAP7_75t_R
XU294 VSS VDD  n340 N138 INVx1_ASAP7_75t_R
XU295 VSS VDD  n342 N139 INVx1_ASAP7_75t_R
XU296 VSS VDD  n343 N140 INVx1_ASAP7_75t_R
XU297 VSS VDD  n339 n344 INVx1_ASAP7_75t_R
XU298 VSS VDD  n341 n345 INVx1_ASAP7_75t_R
XU299 VSS VDD  n346 N74 INVx1_ASAP7_75t_R
XU300 VSS VDD  n348 N75 INVx1_ASAP7_75t_R
XU301 VSS VDD  n350 N76 INVx1_ASAP7_75t_R
XU302 VSS VDD  n351 N77 INVx1_ASAP7_75t_R
XU303 VSS VDD  n347 n352 INVx1_ASAP7_75t_R
XU304 VSS VDD  n349 n353 INVx1_ASAP7_75t_R
XU305 VSS VDD  n354 add_5_root_add_0_root_add_96_31_B_1_ INVx1_ASAP7_75t_R
XU306 VSS VDD  n356 add_5_root_add_0_root_add_96_31_B_2_ INVx1_ASAP7_75t_R
XU307 VSS VDD  n358 add_5_root_add_0_root_add_96_31_B_3_ INVx1_ASAP7_75t_R
XU308 VSS VDD  n360 add_5_root_add_0_root_add_96_31_B_4_ INVx1_ASAP7_75t_R
XU309 VSS VDD  n361 add_5_root_add_0_root_add_96_31_B_5_ INVx1_ASAP7_75t_R
XU310 VSS VDD  n355 n362 INVx1_ASAP7_75t_R
XU311 VSS VDD  n357 n363 INVx1_ASAP7_75t_R
XU312 VSS VDD  n359 n364 INVx1_ASAP7_75t_R
XU313 VSS VDD  n365 add_1_root_add_0_root_add_96_31_B_1_ INVx1_ASAP7_75t_R
XU314 VSS VDD  n367 add_1_root_add_0_root_add_96_31_B_2_ INVx1_ASAP7_75t_R
XU315 VSS VDD  n369 add_1_root_add_0_root_add_96_31_B_3_ INVx1_ASAP7_75t_R
XU316 VSS VDD  n371 add_1_root_add_0_root_add_96_31_B_4_ INVx1_ASAP7_75t_R
XU317 VSS VDD  n373 add_1_root_add_0_root_add_96_31_B_5_ INVx1_ASAP7_75t_R
XU318 VSS VDD  n374 add_1_root_add_0_root_add_96_31_B_6_ INVx1_ASAP7_75t_R
XU319 VSS VDD  n366 n375 INVx1_ASAP7_75t_R
XU320 VSS VDD  n368 n376 INVx1_ASAP7_75t_R
XU321 VSS VDD  n370 n377 INVx1_ASAP7_75t_R
XU322 VSS VDD  n372 n378 INVx1_ASAP7_75t_R
XU323 VSS VDD  n379 N209 INVx1_ASAP7_75t_R
XU324 VSS VDD  n381 N210 INVx1_ASAP7_75t_R
XU325 VSS VDD  n383 N211 INVx1_ASAP7_75t_R
XU326 VSS VDD  n384 N212 INVx1_ASAP7_75t_R
XU327 VSS VDD  n380 n385 INVx1_ASAP7_75t_R
XU328 VSS VDD  n382 n386 INVx1_ASAP7_75t_R
XU329 VSS VDD  n387 N119 INVx1_ASAP7_75t_R
XU330 VSS VDD  n389 N120 INVx1_ASAP7_75t_R
XU331 VSS VDD  n391 N121 INVx1_ASAP7_75t_R
XU332 VSS VDD  n392 N122 INVx1_ASAP7_75t_R
XU333 VSS VDD  n388 n393 INVx1_ASAP7_75t_R
XU334 VSS VDD  n390 n394 INVx1_ASAP7_75t_R
XU335 VSS VDD  n395 add_6_root_add_0_root_add_96_31_B_1_ INVx1_ASAP7_75t_R
XU336 VSS VDD  n397 add_6_root_add_0_root_add_96_31_B_2_ INVx1_ASAP7_75t_R
XU337 VSS VDD  n399 add_6_root_add_0_root_add_96_31_B_3_ INVx1_ASAP7_75t_R
XU338 VSS VDD  n401 add_6_root_add_0_root_add_96_31_B_4_ INVx1_ASAP7_75t_R
XU339 VSS VDD  n402 add_6_root_add_0_root_add_96_31_B_5_ INVx1_ASAP7_75t_R
XU340 VSS VDD  n396 n403 INVx1_ASAP7_75t_R
XU341 VSS VDD  n398 n404 INVx1_ASAP7_75t_R
XU342 VSS VDD  n400 n405 INVx1_ASAP7_75t_R
XU343 VSS VDD  n406 N110 INVx1_ASAP7_75t_R
XU344 VSS VDD  n408 N111 INVx1_ASAP7_75t_R
XU345 VSS VDD  n410 N112 INVx1_ASAP7_75t_R
XU346 VSS VDD  n411 N113 INVx1_ASAP7_75t_R
XU347 VSS VDD  n407 n412 INVx1_ASAP7_75t_R
XU348 VSS VDD  n409 n413 INVx1_ASAP7_75t_R
XU349 VSS VDD  n414 N182 INVx1_ASAP7_75t_R
XU350 VSS VDD  n416 N183 INVx1_ASAP7_75t_R
XU351 VSS VDD  n418 N184 INVx1_ASAP7_75t_R
XU352 VSS VDD  n419 N185 INVx1_ASAP7_75t_R
XU353 VSS VDD  n415 n420 INVx1_ASAP7_75t_R
XU354 VSS VDD  n417 n421 INVx1_ASAP7_75t_R
XU355 VSS VDD  n422 N38 INVx1_ASAP7_75t_R
XU356 VSS VDD  n424 N39 INVx1_ASAP7_75t_R
XU357 VSS VDD  n426 N40 INVx1_ASAP7_75t_R
XU358 VSS VDD  n428 N41 INVx1_ASAP7_75t_R
XU359 VSS VDD  n429 N42 INVx1_ASAP7_75t_R
XU360 VSS VDD  n423 n430 INVx1_ASAP7_75t_R
XU361 VSS VDD  n425 n431 INVx1_ASAP7_75t_R
XU362 VSS VDD  n427 n432 INVx1_ASAP7_75t_R
XU363 VSS VDD  n433 N200 INVx1_ASAP7_75t_R
XU364 VSS VDD  n435 N201 INVx1_ASAP7_75t_R
XU365 VSS VDD  n437 N202 INVx1_ASAP7_75t_R
XU366 VSS VDD  n438 N203 INVx1_ASAP7_75t_R
XU367 VSS VDD  n434 n439 INVx1_ASAP7_75t_R
XU368 VSS VDD  n436 n440 INVx1_ASAP7_75t_R
XU369 VSS VDD  n441 N236 INVx1_ASAP7_75t_R
XU370 VSS VDD  n443 N237 INVx1_ASAP7_75t_R
XU371 VSS VDD  n445 N238 INVx1_ASAP7_75t_R
XU372 VSS VDD  n446 N239 INVx1_ASAP7_75t_R
XU373 VSS VDD  n442 n447 INVx1_ASAP7_75t_R
XU374 VSS VDD  n444 n448 INVx1_ASAP7_75t_R
XU375 VSS VDD  n449 N47 INVx1_ASAP7_75t_R
XU376 VSS VDD  n451 N48 INVx1_ASAP7_75t_R
XU377 VSS VDD  n453 N49 INVx1_ASAP7_75t_R
XU378 VSS VDD  n455 N50 INVx1_ASAP7_75t_R
XU379 VSS VDD  n456 N51 INVx1_ASAP7_75t_R
XU380 VSS VDD  n450 n457 INVx1_ASAP7_75t_R
XU381 VSS VDD  n452 n458 INVx1_ASAP7_75t_R
XU382 VSS VDD  n454 n459 INVx1_ASAP7_75t_R
XU383 VSS VDD  n460 N128 INVx1_ASAP7_75t_R
XU384 VSS VDD  n462 N129 INVx1_ASAP7_75t_R
XU385 VSS VDD  n464 N130 INVx1_ASAP7_75t_R
XU386 VSS VDD  n465 N131 INVx1_ASAP7_75t_R
XU387 VSS VDD  n461 n466 INVx1_ASAP7_75t_R
XU388 VSS VDD  n463 n467 INVx1_ASAP7_75t_R
XU389 VSS VDD  n468 N65 INVx1_ASAP7_75t_R
XU390 VSS VDD  n470 N66 INVx1_ASAP7_75t_R
XU391 VSS VDD  n472 N67 INVx1_ASAP7_75t_R
XU392 VSS VDD  n473 N68 INVx1_ASAP7_75t_R
XU393 VSS VDD  n469 n474 INVx1_ASAP7_75t_R
XU394 VSS VDD  n471 n475 INVx1_ASAP7_75t_R
XU395 VSS VDD  n476 N56 INVx1_ASAP7_75t_R
XU396 VSS VDD  n478 N57 INVx1_ASAP7_75t_R
XU397 VSS VDD  n480 N58 INVx1_ASAP7_75t_R
XU398 VSS VDD  n482 N59 INVx1_ASAP7_75t_R
XU399 VSS VDD  n483 N60 INVx1_ASAP7_75t_R
XU400 VSS VDD  n477 n484 INVx1_ASAP7_75t_R
XU401 VSS VDD  n479 n485 INVx1_ASAP7_75t_R
XU402 VSS VDD  n481 n486 INVx1_ASAP7_75t_R
XU403 VSS VDD  n487 N146 INVx1_ASAP7_75t_R
XU404 VSS VDD  n489 N147 INVx1_ASAP7_75t_R
XU405 VSS VDD  n491 N148 INVx1_ASAP7_75t_R
XU406 VSS VDD  n493 N149 INVx1_ASAP7_75t_R
XU407 VSS VDD  n495 N150 INVx1_ASAP7_75t_R
XU408 VSS VDD  n496 N151 INVx1_ASAP7_75t_R
XU409 VSS VDD  n488 n497 INVx1_ASAP7_75t_R
XU410 VSS VDD  n490 n498 INVx1_ASAP7_75t_R
XU411 VSS VDD  n492 n499 INVx1_ASAP7_75t_R
XU412 VSS VDD  n494 n500 INVx1_ASAP7_75t_R
XU413 VSS VDD  n501 N155 INVx1_ASAP7_75t_R
XU414 VSS VDD  n503 N156 INVx1_ASAP7_75t_R
XU415 VSS VDD  n505 N157 INVx1_ASAP7_75t_R
XU416 VSS VDD  n507 N158 INVx1_ASAP7_75t_R
XU417 VSS VDD  n509 N159 INVx1_ASAP7_75t_R
XU418 VSS VDD  n510 N160 INVx1_ASAP7_75t_R
XU419 VSS VDD  n502 n511 INVx1_ASAP7_75t_R
XU420 VSS VDD  n504 n512 INVx1_ASAP7_75t_R
XU421 VSS VDD  n506 n513 INVx1_ASAP7_75t_R
XU422 VSS VDD  n508 n514 INVx1_ASAP7_75t_R
XU423 VSS VDD  n515 N218 INVx1_ASAP7_75t_R
XU424 VSS VDD  n517 N219 INVx1_ASAP7_75t_R
XU425 VSS VDD  n519 N220 INVx1_ASAP7_75t_R
XU426 VSS VDD  n521 N221 INVx1_ASAP7_75t_R
XU427 VSS VDD  n523 N222 INVx1_ASAP7_75t_R
XU428 VSS VDD  n525 N223 INVx1_ASAP7_75t_R
XU429 VSS VDD  n526 N224 INVx1_ASAP7_75t_R
XU430 VSS VDD  n516 n527 INVx1_ASAP7_75t_R
XU431 VSS VDD  n518 n528 INVx1_ASAP7_75t_R
XU432 VSS VDD  n520 n529 INVx1_ASAP7_75t_R
XU433 VSS VDD  n522 n530 INVx1_ASAP7_75t_R
XU434 VSS VDD  n524 n531 INVx1_ASAP7_75t_R
XU435 VSS VDD  n532 N254 INVx1_ASAP7_75t_R
XU436 VSS VDD  n534 N255 INVx1_ASAP7_75t_R
XU437 VSS VDD  n536 N256 INVx1_ASAP7_75t_R
XU438 VSS VDD  n538 N257 INVx1_ASAP7_75t_R
XU439 VSS VDD  n540 N258 INVx1_ASAP7_75t_R
XU440 VSS VDD  n542 N259 INVx1_ASAP7_75t_R
XU441 VSS VDD  n543 N260 INVx1_ASAP7_75t_R
XU442 VSS VDD  n533 n544 INVx1_ASAP7_75t_R
XU443 VSS VDD  n535 n545 INVx1_ASAP7_75t_R
XU444 VSS VDD  n537 n546 INVx1_ASAP7_75t_R
XU445 VSS VDD  n539 n547 INVx1_ASAP7_75t_R
XU446 VSS VDD  n541 n548 INVx1_ASAP7_75t_R
XU447 VSS VDD  n588 n562 n598 NAND2xp5_ASAP7_75t_R
XU448 VSS VDD  input_buffer[3] n561 n567 NAND2xp5_ASAP7_75t_R
XU449 VSS VDD  input_buffer[4] cnt[0] n566 NAND2xp5_ASAP7_75t_R
XU450 VSS VDD  n567 n566 n600 NAND2xp5_ASAP7_75t_R
XU451 VSS VDD  n600 N6 n571 NAND2xp5_ASAP7_75t_R
XU452 VSS VDD  input_buffer[5] n561 n569 NAND2xp5_ASAP7_75t_R
XU453 VSS VDD  input_buffer[6] cnt[0] n568 NAND2xp5_ASAP7_75t_R
XU454 VSS VDD  n569 n568 n621 NAND2xp5_ASAP7_75t_R
XU455 VSS VDD  n621 n562 n570 NAND2xp5_ASAP7_75t_R
XU456 VSS VDD  n571 n570 n612 NAND2xp5_ASAP7_75t_R
XU457 VSS VDD  input_buffer[7] n561 n573 NAND2xp5_ASAP7_75t_R
XU458 VSS VDD  input_buffer[8] cnt[0] n572 NAND2xp5_ASAP7_75t_R
XU459 VSS VDD  n573 n572 n620 NAND2xp5_ASAP7_75t_R
XU460 VSS VDD  input_buffer[4] n561 n578 NAND2xp5_ASAP7_75t_R
XU461 VSS VDD  input_buffer[5] cnt[0] n577 NAND2xp5_ASAP7_75t_R
XU462 VSS VDD  n578 n577 n607 NAND2xp5_ASAP7_75t_R
XU463 VSS VDD  n607 N6 n582 NAND2xp5_ASAP7_75t_R
XU464 VSS VDD  input_buffer[6] n561 n580 NAND2xp5_ASAP7_75t_R
XU465 VSS VDD  input_buffer[7] cnt[0] n579 NAND2xp5_ASAP7_75t_R
XU466 VSS VDD  n580 n579 n630 NAND2xp5_ASAP7_75t_R
XU467 VSS VDD  n630 n562 n581 NAND2xp5_ASAP7_75t_R
XU468 VSS VDD  n582 n581 n616 NAND2xp5_ASAP7_75t_R
XU469 VSS VDD  input_buffer[8] n561 n629 NAND2xp5_ASAP7_75t_R
XU470 VSS VDD  input_buffer[0] n561 n587 NAND2xp5_ASAP7_75t_R
XU471 VSS VDD  input_buffer[1] cnt[0] n586 NAND2xp5_ASAP7_75t_R
XU472 VSS VDD  n587 n586 n593 NAND2xp5_ASAP7_75t_R
XU473 VSS VDD  n593 n562 n605 NAND2xp5_ASAP7_75t_R
XU474 VSS VDD  n588 N6 n592 NAND2xp5_ASAP7_75t_R
XU475 VSS VDD  input_buffer[1] n561 n590 NAND2xp5_ASAP7_75t_R
XU476 VSS VDD  input_buffer[2] cnt[0] n589 NAND2xp5_ASAP7_75t_R
XU477 VSS VDD  n590 n589 n599 NAND2xp5_ASAP7_75t_R
XU478 VSS VDD  n599 n562 n591 NAND2xp5_ASAP7_75t_R
XU479 VSS VDD  n592 n591 n613 NAND2xp5_ASAP7_75t_R
XU480 VSS VDD  n593 N6 n597 NAND2xp5_ASAP7_75t_R
XU481 VSS VDD  input_buffer[2] n561 n595 NAND2xp5_ASAP7_75t_R
XU482 VSS VDD  input_buffer[3] cnt[0] n594 NAND2xp5_ASAP7_75t_R
XU483 VSS VDD  n595 n594 n606 NAND2xp5_ASAP7_75t_R
XU484 VSS VDD  n606 n562 n596 NAND2xp5_ASAP7_75t_R
XU485 VSS VDD  n597 n596 n617 NAND2xp5_ASAP7_75t_R
XU486 VSS VDD  n599 N6 n602 NAND2xp5_ASAP7_75t_R
XU487 VSS VDD  n600 n562 n601 NAND2xp5_ASAP7_75t_R
XU488 VSS VDD  n602 n601 n625 NAND2xp5_ASAP7_75t_R
XU489 VSS VDD  n606 N6 n609 NAND2xp5_ASAP7_75t_R
XU490 VSS VDD  n607 n562 n608 NAND2xp5_ASAP7_75t_R
XU491 VSS VDD  n609 n608 n628 NAND2xp5_ASAP7_75t_R
XU492 VSS VDD  N279 n549 INVx1_ASAP7_75t_R
XU493 VSS VDD  N278 n550 INVx1_ASAP7_75t_R
XU494 VSS VDD  N277 n551 INVx1_ASAP7_75t_R
XU495 VSS VDD  N276 n552 INVx1_ASAP7_75t_R
XU496 VSS VDD  N275 n553 INVx1_ASAP7_75t_R
XU497 VSS VDD  N274 n554 INVx1_ASAP7_75t_R
XU498 VSS VDD  N273 n555 INVx1_ASAP7_75t_R
XU499 VSS VDD  N272 n556 INVx1_ASAP7_75t_R
XU500 VSS VDD  N271 n557 INVx1_ASAP7_75t_R
XU501 VSS VDD  rst_n n558 INVx1_ASAP7_75t_R
XU502 VSS VDD  n617 n559 INVx1_ASAP7_75t_R
XU503 VSS VDD  n613 n560 INVx1_ASAP7_75t_R
XU504 VSS VDD  n242 n563 INVx1_ASAP7_75t_R
XU505 VSS VDD  n241 n564 INVx1_ASAP7_75t_R
XU506 VSS VDD  n151 n565 INVx1_ASAP7_75t_R
XU507 VSS VDD  input_buffer[0] cnt[0] n588 AND2x2_ASAP7_75t_R
XU508 VSS VDD  n620 N6 n574 AND2x2_ASAP7_75t_R
XU509 VSS VDD  n598 n242 n604 AND2x2_ASAP7_75t_R
XU510 VSS VDD  n605 n242 n611 AND2x2_ASAP7_75t_R
XU511 VSS VDD  n562 n629 n632 AND2x2_ASAP7_75t_R
.ENDS


.SUBCKT VSS VDD  CIM_adder_tree_DW01_add_1 A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] CO
XU1_7 VSS VDD  A[7] B[7] n3 n9 n10 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] n4 n11 n12 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] n5 n13 n14 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] n6 n15 n16 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] n7 n17 n18 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] n8 n19 n20 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] n1 n21 n22 FAx1_ASAP7_75t_R
XU1 VSS VDD  A[0] B[0] n1 AND2x2_ASAP7_75t_R
XU2 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU3 VSS VDD  n11 n3 INVx1_ASAP7_75t_R
XU4 VSS VDD  n13 n4 INVx1_ASAP7_75t_R
XU5 VSS VDD  n15 n5 INVx1_ASAP7_75t_R
XU6 VSS VDD  n17 n6 INVx1_ASAP7_75t_R
XU7 VSS VDD  n19 n7 INVx1_ASAP7_75t_R
XU8 VSS VDD  n21 n8 INVx1_ASAP7_75t_R
XU9 VSS VDD  n9 SUM[8] INVx1_ASAP7_75t_R
XU10 VSS VDD  n10 SUM[7] INVx1_ASAP7_75t_R
XU11 VSS VDD  n12 SUM[6] INVx1_ASAP7_75t_R
XU12 VSS VDD  n14 SUM[5] INVx1_ASAP7_75t_R
XU13 VSS VDD  n16 SUM[4] INVx1_ASAP7_75t_R
XU14 VSS VDD  n18 SUM[3] INVx1_ASAP7_75t_R
XU15 VSS VDD  n20 SUM[2] INVx1_ASAP7_75t_R
XU16 VSS VDD  n22 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT VSS VDD  CIM_adder_tree_DW01_add_0 A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[12] SUM[11] SUM[10] SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] CO
XU1_11 VSS VDD  A[11] B[11] n5 n15 n16 FAx1_ASAP7_75t_R
XU1_10 VSS VDD  A[10] B[10] n6 n17 n18 FAx1_ASAP7_75t_R
XU1_9 VSS VDD  A[9] B[9] n7 n19 n20 FAx1_ASAP7_75t_R
XU1_8 VSS VDD  A[8] B[8] n8 n21 n22 FAx1_ASAP7_75t_R
XU1_7 VSS VDD  A[7] B[7] n9 n23 n24 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] n10 n25 n26 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] n11 n27 n28 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] n12 n29 n30 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] n13 n31 n32 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] n14 n33 n34 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] n1 n35 n36 FAx1_ASAP7_75t_R
XU1 VSS VDD  A[0] B[0] n1 AND2x2_ASAP7_75t_R
XU2 VSS VDD  A[12] n4 SUM[12] XOR2xp5_ASAP7_75t_R
XU3 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU4 VSS VDD  n15 n4 INVx1_ASAP7_75t_R
XU5 VSS VDD  n17 n5 INVx1_ASAP7_75t_R
XU6 VSS VDD  n19 n6 INVx1_ASAP7_75t_R
XU7 VSS VDD  n21 n7 INVx1_ASAP7_75t_R
XU8 VSS VDD  n23 n8 INVx1_ASAP7_75t_R
XU9 VSS VDD  n25 n9 INVx1_ASAP7_75t_R
XU10 VSS VDD  n27 n10 INVx1_ASAP7_75t_R
XU11 VSS VDD  n29 n11 INVx1_ASAP7_75t_R
XU12 VSS VDD  n31 n12 INVx1_ASAP7_75t_R
XU13 VSS VDD  n33 n13 INVx1_ASAP7_75t_R
XU14 VSS VDD  n35 n14 INVx1_ASAP7_75t_R
XU15 VSS VDD  n20 SUM[9] INVx1_ASAP7_75t_R
XU16 VSS VDD  n22 SUM[8] INVx1_ASAP7_75t_R
XU17 VSS VDD  n24 SUM[7] INVx1_ASAP7_75t_R
XU18 VSS VDD  n26 SUM[6] INVx1_ASAP7_75t_R
XU19 VSS VDD  n28 SUM[5] INVx1_ASAP7_75t_R
XU20 VSS VDD  n30 SUM[4] INVx1_ASAP7_75t_R
XU21 VSS VDD  n32 SUM[3] INVx1_ASAP7_75t_R
XU22 VSS VDD  n34 SUM[2] INVx1_ASAP7_75t_R
XU23 VSS VDD  n36 SUM[1] INVx1_ASAP7_75t_R
XU24 VSS VDD  n16 SUM[11] INVx1_ASAP7_75t_R
XU25 VSS VDD  n18 SUM[10] INVx1_ASAP7_75t_R
.ENDS


