.SUBCKT CIM_adder_tree rst_n clk Input_1[3] Input_1[2] Input_1[1] Input_1[0] Input_2[3] Input_2[2] Input_2[1] Input_2[0] Input_3[3] Input_3[2] Input_3[1] Input_3[0] Input_4[3] Input_4[2] Input_4[1] Input_4[0] Input_5[3] Input_5[2] Input_5[1] Input_5[0] Input_6[3] Input_6[2] Input_6[1] Input_6[0] Input_7[3] Input_7[2] Input_7[1] Input_7[0] Input_8[3] Input_8[2] Input_8[1] Input_8[0] Input_9[3] Input_9[2] Input_9[1] Input_9[0] Input_10[3] Input_10[2] Input_10[1] Input_10[0] Input_11[3] Input_11[2] Input_11[1] Input_11[0] Input_12[3] Input_12[2] Input_12[1] Input_12[0] Input_13[3] Input_13[2] Input_13[1] Input_13[0] Input_14[3] Input_14[2] Input_14[1] Input_14[0] Input_15[3] Input_15[2] Input_15[1] Input_15[0] Input_16[3] Input_16[2] Input_16[1] Input_16[0] Input_17[3] Input_17[2] Input_17[1] Input_17[0] Input_18[3] Input_18[2] Input_18[1] Input_18[0] Input_19[3] Input_19[2] Input_19[1] Input_19[0] Input_20[3] Input_20[2] Input_20[1] Input_20[0] Input_21[3] Input_21[2] Input_21[1] Input_21[0] Input_22[3] Input_22[2] Input_22[1] Input_22[0] Input_23[3] Input_23[2] Input_23[1] Input_23[0] Input_24[3] Input_24[2] Input_24[1] Input_24[0] Input_25[3] Input_25[2] Input_25[1] Input_25[0] Input_26[3] Input_26[2] Input_26[1] Input_26[0] Input_27[3] Input_27[2] Input_27[1] Input_27[0] Input_28[3] Input_28[2] Input_28[1] Input_28[0] Input_29[3] Input_29[2] Input_29[1] Input_29[0] Input_30[3] Input_30[2] Input_30[1] Input_30[0] Input_31[3] Input_31[2] Input_31[1] Input_31[0] Input_32[3] Input_32[2] Input_32[1] Input_32[0] out_valid Output[12] Output[11] Output[10] Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0]
XU82 cnt[1] cnt[0] n149 NAND2xp5_ASAP7_75t_R
XU85 cnt[2] n565 n152 NAND2xp5_ASAP7_75t_R
Xadd_123 Output[12] Output[11] Output[10] Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0] n233 shift_buffer[11] shift_buffer[10] shift_buffer[9] shift_buffer[8] shift_buffer[7] shift_buffer[6] shift_buffer[5] shift_buffer[4] shift_buffer[3] shift_buffer[2] shift_buffer[1] shift_buffer[0] n233 N309 N308 N307 N306 N305 N304 N303 N302 N301 N300 N299 N298 N297 CIM_adder_tree_DW01_add_0
Xadd_0_root_add_0_root_add_96_31 n233 N224 N223 N222 N221 N220 N219 N218 n167 n233 N260 N259 N258 N257 N256 N255 N254 n182 n233 N279 N278 N277 N276 N275 N274 N273 N272 N271 CIM_adder_tree_DW01_add_1
Xadd_1_root_add_0_root_add_96_31_U1_1 add_1_root_add_0_root_add_96_31_A_1_ add_1_root_add_0_root_add_96_31_B_1_ n165 n533 n532 FAx1_ASAP7_75t_R
Xadd_1_root_add_0_root_add_96_31_U1_2 add_1_root_add_0_root_add_96_31_A_2_ add_1_root_add_0_root_add_96_31_B_2_ n544 n535 n534 FAx1_ASAP7_75t_R
Xadd_1_root_add_0_root_add_96_31_U1_3 add_1_root_add_0_root_add_96_31_A_3_ add_1_root_add_0_root_add_96_31_B_3_ n545 n537 n536 FAx1_ASAP7_75t_R
Xadd_1_root_add_0_root_add_96_31_U1_4 add_1_root_add_0_root_add_96_31_A_4_ add_1_root_add_0_root_add_96_31_B_4_ n546 n539 n538 FAx1_ASAP7_75t_R
Xadd_1_root_add_0_root_add_96_31_U1_5 add_1_root_add_0_root_add_96_31_A_5_ add_1_root_add_0_root_add_96_31_B_5_ n547 n541 n540 FAx1_ASAP7_75t_R
Xadd_1_root_add_0_root_add_96_31_U1_6 add_1_root_add_0_root_add_96_31_A_6_ add_1_root_add_0_root_add_96_31_B_6_ n548 n543 n542 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_1 N155 N146 n166 n516 n515 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_2 N156 N147 n527 n518 n517 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_3 N157 N148 n528 n520 n519 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_4 N158 N149 n529 n522 n521 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_5 N159 N150 n530 n524 n523 FAx1_ASAP7_75t_R
Xadd_2_root_add_0_root_add_96_31_U1_6 N160 N151 n531 n526 n525 FAx1_ASAP7_75t_R
Xadd_6_root_add_0_root_add_96_31_U1_1 N47 add_6_root_add_0_root_add_96_31_B_1_ n164 n502 n501 FAx1_ASAP7_75t_R
Xadd_6_root_add_0_root_add_96_31_U1_2 N48 add_6_root_add_0_root_add_96_31_B_2_ n511 n504 n503 FAx1_ASAP7_75t_R
Xadd_6_root_add_0_root_add_96_31_U1_3 N49 add_6_root_add_0_root_add_96_31_B_3_ n512 n506 n505 FAx1_ASAP7_75t_R
Xadd_6_root_add_0_root_add_96_31_U1_4 N50 add_6_root_add_0_root_add_96_31_B_4_ n513 n508 n507 FAx1_ASAP7_75t_R
Xadd_6_root_add_0_root_add_96_31_U1_5 N51 add_6_root_add_0_root_add_96_31_B_5_ n514 n510 n509 FAx1_ASAP7_75t_R
Xadd_3_root_add_0_root_add_96_31_U1_1 N56 N38 n163 n488 n487 FAx1_ASAP7_75t_R
Xadd_3_root_add_0_root_add_96_31_U1_2 N57 N39 n497 n490 n489 FAx1_ASAP7_75t_R
Xadd_3_root_add_0_root_add_96_31_U1_3 N58 N40 n498 n492 n491 FAx1_ASAP7_75t_R
Xadd_3_root_add_0_root_add_96_31_U1_4 N59 N41 n499 n494 n493 FAx1_ASAP7_75t_R
Xadd_3_root_add_0_root_add_96_31_U1_5 N60 N42 n500 n496 n495 FAx1_ASAP7_75t_R
Xadd_14_root_add_0_root_add_96_31_U1_1 N128 N65 n158 n477 n476 FAx1_ASAP7_75t_R
Xadd_14_root_add_0_root_add_96_31_U1_2 N129 N66 n484 n479 n478 FAx1_ASAP7_75t_R
Xadd_14_root_add_0_root_add_96_31_U1_3 N130 N67 n485 n481 n480 FAx1_ASAP7_75t_R
Xadd_14_root_add_0_root_add_96_31_U1_4 N131 N68 n486 n483 n482 FAx1_ASAP7_75t_R
Xadd_15_root_add_0_root_add_96_31_U1_1 Input_15[1] Input_14[1] n197 n469 n468 FAx1_ASAP7_75t_R
Xadd_15_root_add_0_root_add_96_31_U1_2 Input_15[2] Input_14[2] n474 n471 n470 FAx1_ASAP7_75t_R
Xadd_15_root_add_0_root_add_96_31_U1_3 Input_15[3] Input_14[3] n475 n473 n472 FAx1_ASAP7_75t_R
Xadd_29_root_add_0_root_add_96_31_U1_1 Input_30[1] Input_2[1] n193 n461 n460 FAx1_ASAP7_75t_R
Xadd_29_root_add_0_root_add_96_31_U1_2 Input_30[2] Input_2[2] n466 n463 n462 FAx1_ASAP7_75t_R
Xadd_29_root_add_0_root_add_96_31_U1_3 Input_30[3] Input_2[3] n467 n465 n464 FAx1_ASAP7_75t_R
Xadd_12_root_add_0_root_add_96_31_U1_1 N200 N236 n157 n450 n449 FAx1_ASAP7_75t_R
Xadd_12_root_add_0_root_add_96_31_U1_2 N201 N237 n457 n452 n451 FAx1_ASAP7_75t_R
Xadd_12_root_add_0_root_add_96_31_U1_3 N202 N238 n458 n454 n453 FAx1_ASAP7_75t_R
Xadd_12_root_add_0_root_add_96_31_U1_4 N203 N239 n459 n456 n455 FAx1_ASAP7_75t_R
Xadd_17_root_add_0_root_add_96_31_U1_1 Input_12[1] Input_6[1] n196 n442 n441 FAx1_ASAP7_75t_R
Xadd_17_root_add_0_root_add_96_31_U1_2 Input_12[2] Input_6[2] n447 n444 n443 FAx1_ASAP7_75t_R
Xadd_17_root_add_0_root_add_96_31_U1_3 Input_12[3] Input_6[3] n448 n446 n445 FAx1_ASAP7_75t_R
Xadd_25_root_add_0_root_add_96_31_U1_1 Input_26[1] Input_17[1] n192 n434 n433 FAx1_ASAP7_75t_R
Xadd_25_root_add_0_root_add_96_31_U1_2 Input_26[2] Input_17[2] n439 n436 n435 FAx1_ASAP7_75t_R
Xadd_25_root_add_0_root_add_96_31_U1_3 Input_26[3] Input_17[3] n440 n438 n437 FAx1_ASAP7_75t_R
Xadd_11_root_add_0_root_add_96_31_U1_1 N110 N182 n160 n423 n422 FAx1_ASAP7_75t_R
Xadd_11_root_add_0_root_add_96_31_U1_2 N111 N183 n430 n425 n424 FAx1_ASAP7_75t_R
Xadd_11_root_add_0_root_add_96_31_U1_3 N112 N184 n431 n427 n426 FAx1_ASAP7_75t_R
Xadd_11_root_add_0_root_add_96_31_U1_4 N113 N185 n432 n429 n428 FAx1_ASAP7_75t_R
Xadd_18_root_add_0_root_add_96_31_U1_1 Input_3[1] Input_21[1] n199 n415 n414 FAx1_ASAP7_75t_R
Xadd_18_root_add_0_root_add_96_31_U1_2 Input_3[2] Input_21[2] n420 n417 n416 FAx1_ASAP7_75t_R
Xadd_18_root_add_0_root_add_96_31_U1_3 Input_3[3] Input_21[3] n421 n419 n418 FAx1_ASAP7_75t_R
Xadd_26_root_add_0_root_add_96_31_U1_1 Input_27[1] Input_16[1] n195 n407 n406 FAx1_ASAP7_75t_R
Xadd_26_root_add_0_root_add_96_31_U1_2 Input_27[2] Input_16[2] n412 n409 n408 FAx1_ASAP7_75t_R
Xadd_26_root_add_0_root_add_96_31_U1_3 Input_27[3] Input_16[3] n413 n411 n410 FAx1_ASAP7_75t_R
Xadd_7_root_add_0_root_add_96_31_U1_1 N209 N119 n159 n396 n395 FAx1_ASAP7_75t_R
Xadd_7_root_add_0_root_add_96_31_U1_2 N210 N120 n403 n398 n397 FAx1_ASAP7_75t_R
Xadd_7_root_add_0_root_add_96_31_U1_3 N211 N121 n404 n400 n399 FAx1_ASAP7_75t_R
Xadd_7_root_add_0_root_add_96_31_U1_4 N212 N122 n405 n402 n401 FAx1_ASAP7_75t_R
Xadd_27_root_add_0_root_add_96_31_U1_1 Input_28[1] Input_8[1] n198 n388 n387 FAx1_ASAP7_75t_R
Xadd_27_root_add_0_root_add_96_31_U1_2 Input_28[2] Input_8[2] n393 n390 n389 FAx1_ASAP7_75t_R
Xadd_27_root_add_0_root_add_96_31_U1_3 Input_28[3] Input_8[3] n394 n392 n391 FAx1_ASAP7_75t_R
Xadd_28_root_add_0_root_add_96_31_U1_1 Input_29[1] Input_4[1] n194 n380 n379 FAx1_ASAP7_75t_R
Xadd_28_root_add_0_root_add_96_31_U1_2 Input_29[2] Input_4[2] n385 n382 n381 FAx1_ASAP7_75t_R
Xadd_28_root_add_0_root_add_96_31_U1_3 Input_29[3] Input_4[3] n386 n384 n383 FAx1_ASAP7_75t_R
Xadd_5_root_add_0_root_add_96_31_U1_1 N173 add_5_root_add_0_root_add_96_31_B_1_ n161 n366 n365 FAx1_ASAP7_75t_R
Xadd_5_root_add_0_root_add_96_31_U1_2 N174 add_5_root_add_0_root_add_96_31_B_2_ n375 n368 n367 FAx1_ASAP7_75t_R
Xadd_5_root_add_0_root_add_96_31_U1_3 N175 add_5_root_add_0_root_add_96_31_B_3_ n376 n370 n369 FAx1_ASAP7_75t_R
Xadd_5_root_add_0_root_add_96_31_U1_4 N176 add_5_root_add_0_root_add_96_31_B_4_ n377 n372 n371 FAx1_ASAP7_75t_R
Xadd_5_root_add_0_root_add_96_31_U1_5 N177 add_5_root_add_0_root_add_96_31_B_5_ n378 n374 n373 FAx1_ASAP7_75t_R
Xadd_8_root_add_0_root_add_96_31_U1_1 N137 N74 n156 n355 n354 FAx1_ASAP7_75t_R
Xadd_8_root_add_0_root_add_96_31_U1_2 N138 N75 n362 n357 n356 FAx1_ASAP7_75t_R
Xadd_8_root_add_0_root_add_96_31_U1_3 N139 N76 n363 n359 n358 FAx1_ASAP7_75t_R
Xadd_8_root_add_0_root_add_96_31_U1_4 N140 N77 n364 n361 n360 FAx1_ASAP7_75t_R
Xadd_19_root_add_0_root_add_96_31_U1_1 Input_31[1] Input_11[1] n191 n347 n346 FAx1_ASAP7_75t_R
Xadd_19_root_add_0_root_add_96_31_U1_2 Input_31[2] Input_11[2] n352 n349 n348 FAx1_ASAP7_75t_R
Xadd_19_root_add_0_root_add_96_31_U1_3 Input_31[3] Input_11[3] n353 n351 n350 FAx1_ASAP7_75t_R
Xadd_30_root_add_0_root_add_96_31_U1_1 Input_1[1] Input_32[1] n187 n339 n338 FAx1_ASAP7_75t_R
Xadd_30_root_add_0_root_add_96_31_U1_2 Input_1[2] Input_32[2] n344 n341 n340 FAx1_ASAP7_75t_R
Xadd_30_root_add_0_root_add_96_31_U1_3 Input_1[3] Input_32[3] n345 n343 n342 FAx1_ASAP7_75t_R
Xadd_13_root_add_0_root_add_96_31_U1_1 N245 N263 n154 n328 n327 FAx1_ASAP7_75t_R
Xadd_13_root_add_0_root_add_96_31_U1_2 N246 N264 n335 n330 n329 FAx1_ASAP7_75t_R
Xadd_13_root_add_0_root_add_96_31_U1_3 N247 N265 n336 n332 n331 FAx1_ASAP7_75t_R
Xadd_13_root_add_0_root_add_96_31_U1_4 N248 N266 n337 n334 n333 FAx1_ASAP7_75t_R
Xadd_16_root_add_0_root_add_96_31_U1_1 Input_7[1] Input_13[1] n189 n320 n319 FAx1_ASAP7_75t_R
Xadd_16_root_add_0_root_add_96_31_U1_2 Input_7[2] Input_13[2] n325 n322 n321 FAx1_ASAP7_75t_R
Xadd_16_root_add_0_root_add_96_31_U1_3 Input_7[3] Input_13[3] n326 n324 n323 FAx1_ASAP7_75t_R
Xadd_24_root_add_0_root_add_96_31_U1_1 Input_25[1] Input_9[1] n185 n312 n311 FAx1_ASAP7_75t_R
Xadd_24_root_add_0_root_add_96_31_U1_2 Input_25[2] Input_9[2] n317 n314 n313 FAx1_ASAP7_75t_R
Xadd_24_root_add_0_root_add_96_31_U1_3 Input_25[3] Input_9[3] n318 n316 n315 FAx1_ASAP7_75t_R
Xadd_4_root_add_0_root_add_96_31_U1_1 N164 N227 n162 n298 n297 FAx1_ASAP7_75t_R
Xadd_4_root_add_0_root_add_96_31_U1_2 N165 N228 n307 n300 n299 FAx1_ASAP7_75t_R
Xadd_4_root_add_0_root_add_96_31_U1_3 N166 N229 n308 n302 n301 FAx1_ASAP7_75t_R
Xadd_4_root_add_0_root_add_96_31_U1_4 N167 N230 n309 n304 n303 FAx1_ASAP7_75t_R
Xadd_4_root_add_0_root_add_96_31_U1_5 N168 N231 n310 n306 n305 FAx1_ASAP7_75t_R
Xadd_9_root_add_0_root_add_96_31_U1_1 N83 N101 n155 n287 n286 FAx1_ASAP7_75t_R
Xadd_9_root_add_0_root_add_96_31_U1_2 N84 N102 n294 n289 n288 FAx1_ASAP7_75t_R
Xadd_9_root_add_0_root_add_96_31_U1_3 N85 N103 n295 n291 n290 FAx1_ASAP7_75t_R
Xadd_9_root_add_0_root_add_96_31_U1_4 N86 N104 n296 n293 n292 FAx1_ASAP7_75t_R
Xadd_23_root_add_0_root_add_96_31_U1_1 Input_24[1] Input_18[1] n190 n279 n278 FAx1_ASAP7_75t_R
Xadd_23_root_add_0_root_add_96_31_U1_2 Input_24[2] Input_18[2] n284 n281 n280 FAx1_ASAP7_75t_R
Xadd_23_root_add_0_root_add_96_31_U1_3 Input_24[3] Input_18[3] n285 n283 n282 FAx1_ASAP7_75t_R
Xadd_20_root_add_0_root_add_96_31_U1_1 Input_10[1] Input_20[1] n186 n271 n270 FAx1_ASAP7_75t_R
Xadd_20_root_add_0_root_add_96_31_U1_2 Input_10[2] Input_20[2] n276 n273 n272 FAx1_ASAP7_75t_R
Xadd_20_root_add_0_root_add_96_31_U1_3 Input_10[3] Input_20[3] n277 n275 n274 FAx1_ASAP7_75t_R
Xadd_10_root_add_0_root_add_96_31_U1_1 N92 N191 n153 n260 n259 FAx1_ASAP7_75t_R
Xadd_10_root_add_0_root_add_96_31_U1_2 N93 N192 n267 n262 n261 FAx1_ASAP7_75t_R
Xadd_10_root_add_0_root_add_96_31_U1_3 N94 N193 n268 n264 n263 FAx1_ASAP7_75t_R
Xadd_10_root_add_0_root_add_96_31_U1_4 N95 N194 n269 n266 n265 FAx1_ASAP7_75t_R
Xadd_21_root_add_0_root_add_96_31_U1_1 Input_22[1] Input_5[1] n188 n252 n251 FAx1_ASAP7_75t_R
Xadd_21_root_add_0_root_add_96_31_U1_2 Input_22[2] Input_5[2] n257 n254 n253 FAx1_ASAP7_75t_R
Xadd_21_root_add_0_root_add_96_31_U1_3 Input_22[3] Input_5[3] n258 n256 n255 FAx1_ASAP7_75t_R
Xadd_22_root_add_0_root_add_96_31_U1_1 Input_23[1] Input_19[1] n184 n244 n243 FAx1_ASAP7_75t_R
Xadd_22_root_add_0_root_add_96_31_U1_2 Input_23[2] Input_19[2] n249 n246 n245 FAx1_ASAP7_75t_R
Xadd_22_root_add_0_root_add_96_31_U1_3 Input_23[3] Input_19[3] n250 n248 n247 FAx1_ASAP7_75t_R
Xcnt_reg_0_ n240 clk n233 n558 cnt[0] ASYNC_DFFHx1_ASAP7_75t_R
Xcnt_reg_2_ n563 clk n233 n558 cnt[2] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_2_ n232 clk n558 n233 Output[2] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_1_ n231 clk n558 n233 Output[1] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_0_ n183 clk n558 n233 Output[0] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_3_ n230 clk n558 n233 Output[3] ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg n564 clk n558 n233 out_valid ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_4_ n228 clk n558 n233 Output[4] ASYNC_DFFHx1_ASAP7_75t_R
Xcnt_reg_1_ n229 clk n558 n233 cnt[1] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_5_ n227 clk n558 n233 Output[5] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_6_ n226 clk n558 n233 Output[6] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_3_ n239 clk n558 n233 shift_buffer[3] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_2_ n238 clk n558 n233 shift_buffer[2] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_1_ n237 clk n558 n233 shift_buffer[1] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_0_ n236 clk n558 n233 shift_buffer[0] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_5_ n235 clk n558 n233 shift_buffer[5] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_4_ n234 clk n558 n233 shift_buffer[4] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_7_ n225 clk n558 n233 Output[7] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_11_ n224 clk n558 n233 shift_buffer[11] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_10_ n223 clk n558 n233 shift_buffer[10] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_9_ n222 clk n558 n233 shift_buffer[9] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_8_ n221 clk n558 n233 shift_buffer[8] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_7_ n220 clk n558 n233 shift_buffer[7] ASYNC_DFFHx1_ASAP7_75t_R
Xshift_buffer_reg_6_ n219 clk n558 n233 shift_buffer[6] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_8_ n218 clk n558 n233 Output[8] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_9_ n217 clk n558 n233 Output[9] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_10_ n216 clk n558 n233 Output[10] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_11_ n215 clk n558 n233 Output[11] ASYNC_DFFHx1_ASAP7_75t_R
XOutput_reg_12_ n214 clk n558 n233 Output[12] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_0_ n557 clk n558 n233 input_buffer[0] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_1_ n556 clk n558 n233 input_buffer[1] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_2_ n555 clk n558 n233 input_buffer[2] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_3_ n554 clk n558 n233 input_buffer[3] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_4_ n553 clk n558 n233 input_buffer[4] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_5_ n552 clk n558 n233 input_buffer[5] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_6_ n551 clk n558 n233 input_buffer[6] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_8_ n549 clk n558 n233 input_buffer[8] ASYNC_DFFHx1_ASAP7_75t_R
Xinput_buffer_reg_7_ n550 clk n558 n233 input_buffer[7] ASYNC_DFFHx1_ASAP7_75t_R
XU106 n233 TIELOx1_ASAP7_75t_R
XU107 n242 n625 n603 NOR2xp33_ASAP7_75t_R
XU108 n242 n628 n610 NOR2xp33_ASAP7_75t_R
XU109 n169 n201 n153 AND2x2_ASAP7_75t_R
XU110 n168 n200 n154 AND2x2_ASAP7_75t_R
XU111 n171 n203 n155 AND2x2_ASAP7_75t_R
XU112 n170 n202 n156 AND2x2_ASAP7_75t_R
XU113 n173 n205 n157 AND2x2_ASAP7_75t_R
XU114 n172 n204 n158 AND2x2_ASAP7_75t_R
XU115 n175 n207 n159 AND2x2_ASAP7_75t_R
XU116 n174 n206 n160 AND2x2_ASAP7_75t_R
XU117 n176 n208 n161 AND2x2_ASAP7_75t_R
XU118 n177 n209 n162 AND2x2_ASAP7_75t_R
XU119 n178 n210 n163 AND2x2_ASAP7_75t_R
XU120 n179 n211 n164 AND2x2_ASAP7_75t_R
XU121 n180 n212 n165 AND2x2_ASAP7_75t_R
XU122 n181 n213 n166 AND2x2_ASAP7_75t_R
XU123 n181 n213 n167 XOR2xp5_ASAP7_75t_R
XU124 Input_25[0] Input_9[0] n168 XOR2xp5_ASAP7_75t_R
XU125 Input_23[0] Input_19[0] n169 XOR2xp5_ASAP7_75t_R
XU126 Input_1[0] Input_32[0] n170 XOR2xp5_ASAP7_75t_R
XU127 Input_10[0] Input_20[0] n171 XOR2xp5_ASAP7_75t_R
XU128 Input_30[0] Input_2[0] n172 XOR2xp5_ASAP7_75t_R
XU129 Input_26[0] Input_17[0] n173 XOR2xp5_ASAP7_75t_R
XU130 Input_27[0] Input_16[0] n174 XOR2xp5_ASAP7_75t_R
XU131 Input_29[0] Input_4[0] n175 XOR2xp5_ASAP7_75t_R
XU132 n168 n200 n176 XOR2xp5_ASAP7_75t_R
XU133 n169 n201 n177 XOR2xp5_ASAP7_75t_R
XU134 n172 n204 n178 XOR2xp5_ASAP7_75t_R
XU135 n173 n205 n179 XOR2xp5_ASAP7_75t_R
XU136 n177 n209 n180 XOR2xp5_ASAP7_75t_R
XU137 n179 n211 n181 XOR2xp5_ASAP7_75t_R
XU138 n180 n212 n182 XOR2xp5_ASAP7_75t_R
XU139 N297 n150 n183 NAND2xp5_ASAP7_75t_R
XU140 Input_23[0] Input_19[0] n184 AND2x2_ASAP7_75t_R
XU141 Input_25[0] Input_9[0] n185 AND2x2_ASAP7_75t_R
XU142 Input_10[0] Input_20[0] n186 AND2x2_ASAP7_75t_R
XU143 Input_1[0] Input_32[0] n187 AND2x2_ASAP7_75t_R
XU144 Input_22[0] Input_5[0] n188 AND2x2_ASAP7_75t_R
XU145 Input_7[0] Input_13[0] n189 AND2x2_ASAP7_75t_R
XU146 Input_24[0] Input_18[0] n190 AND2x2_ASAP7_75t_R
XU147 Input_31[0] Input_11[0] n191 AND2x2_ASAP7_75t_R
XU148 Input_26[0] Input_17[0] n192 AND2x2_ASAP7_75t_R
XU149 Input_30[0] Input_2[0] n193 AND2x2_ASAP7_75t_R
XU150 Input_29[0] Input_4[0] n194 AND2x2_ASAP7_75t_R
XU151 Input_27[0] Input_16[0] n195 AND2x2_ASAP7_75t_R
XU152 Input_12[0] Input_6[0] n196 AND2x2_ASAP7_75t_R
XU153 Input_15[0] Input_14[0] n197 AND2x2_ASAP7_75t_R
XU154 Input_28[0] Input_8[0] n198 AND2x2_ASAP7_75t_R
XU155 Input_3[0] Input_21[0] n199 AND2x2_ASAP7_75t_R
XU156 Input_7[0] Input_13[0] n200 XOR2xp5_ASAP7_75t_R
XU157 Input_22[0] Input_5[0] n201 XOR2xp5_ASAP7_75t_R
XU158 Input_31[0] Input_11[0] n202 XOR2xp5_ASAP7_75t_R
XU159 Input_24[0] Input_18[0] n203 XOR2xp5_ASAP7_75t_R
XU160 Input_15[0] Input_14[0] n204 XOR2xp5_ASAP7_75t_R
XU161 Input_12[0] Input_6[0] n205 XOR2xp5_ASAP7_75t_R
XU162 Input_3[0] Input_21[0] n206 XOR2xp5_ASAP7_75t_R
XU163 Input_28[0] Input_8[0] n207 XOR2xp5_ASAP7_75t_R
XU164 n170 n202 n208 XOR2xp5_ASAP7_75t_R
XU165 n171 n203 n209 XOR2xp5_ASAP7_75t_R
XU166 n174 n206 n210 XOR2xp5_ASAP7_75t_R
XU167 n175 n207 n211 XOR2xp5_ASAP7_75t_R
XU168 n176 n208 n212 XOR2xp5_ASAP7_75t_R
XU169 n178 n210 n213 XOR2xp5_ASAP7_75t_R
XU170 N309 n150 n214 NAND2xp5_ASAP7_75t_R
XU171 N308 n150 n215 NAND2xp5_ASAP7_75t_R
XU172 N307 n150 n216 NAND2xp5_ASAP7_75t_R
XU173 N306 n150 n217 NAND2xp5_ASAP7_75t_R
XU174 N305 n150 n218 NAND2xp5_ASAP7_75t_R
XU175 n241 n615 n614 n219 OR3x1_ASAP7_75t_R
XU176 n241 n619 n618 n220 OR3x1_ASAP7_75t_R
XU177 n241 n627 n626 n221 OR3x1_ASAP7_75t_R
XU178 n241 n635 n634 n222 OR3x1_ASAP7_75t_R
XU179 n241 n576 n575 n223 OR3x1_ASAP7_75t_R
XU180 n241 n585 n584 n224 OR3x1_ASAP7_75t_R
XU181 N304 n150 n225 NAND2xp5_ASAP7_75t_R
XU182 N303 n150 n226 NAND2xp5_ASAP7_75t_R
XU183 N302 n150 n227 NAND2xp5_ASAP7_75t_R
XU184 N301 n150 n228 NAND2xp5_ASAP7_75t_R
XU185 n564 N6 n229 NAND2xp5_ASAP7_75t_R
XU186 N300 n150 n230 NAND2xp5_ASAP7_75t_R
XU187 N298 n150 n231 NAND2xp5_ASAP7_75t_R
XU188 N299 n150 n232 NAND2xp5_ASAP7_75t_R
XU189 n242 n612 n615 NOR2xp33_ASAP7_75t_R
XU190 n613 n563 n614 NOR2xp33_ASAP7_75t_R
XU191 n242 n616 n619 NOR2xp33_ASAP7_75t_R
XU192 n617 n563 n618 NOR2xp33_ASAP7_75t_R
XU193 n242 n624 n627 NOR2xp33_ASAP7_75t_R
XU194 n625 n563 n626 NOR2xp33_ASAP7_75t_R
XU195 n242 n583 n584 NOR2xp33_ASAP7_75t_R
XU196 n616 n563 n585 NOR2xp33_ASAP7_75t_R
XU197 n242 n633 n634 NOR2xp33_ASAP7_75t_R
XU198 n628 n563 n635 NOR2xp33_ASAP7_75t_R
XU199 n242 n574 n575 NOR2xp33_ASAP7_75t_R
XU200 n612 n563 n576 NOR2xp33_ASAP7_75t_R
XU201 n241 n604 n603 n234 OR3x1_ASAP7_75t_R
XU202 n241 n611 n610 n235 OR3x1_ASAP7_75t_R
XU203 n598 n241 n242 n236 OR3x1_ASAP7_75t_R
XU204 n605 n241 n242 n237 OR3x1_ASAP7_75t_R
XU205 n560 n241 n242 n238 OR3x1_ASAP7_75t_R
XU206 n559 n241 n242 n239 OR3x1_ASAP7_75t_R
XU207 N6 n562 INVx1_ASAP7_75t_R
XU208 n632 n631 n633 NOR2xp33_ASAP7_75t_R
XU209 n562 n630 n631 NOR2xp33_ASAP7_75t_R
XU210 n623 n622 n624 NOR2xp33_ASAP7_75t_R
XU211 N6 n620 n623 NOR2xp33_ASAP7_75t_R
XU212 n562 n621 n622 NOR2xp33_ASAP7_75t_R
XU213 n562 n629 n583 NOR2xp33_ASAP7_75t_R
XU214 cnt[1] cnt[0] n151 NOR2xp33_ASAP7_75t_R
XU215 N284 n241 HB1xp67_ASAP7_75t_R
XU216 n565 cnt[2] N284 NOR2xp33_ASAP7_75t_R
XU217 N7 n242 HB1xp67_ASAP7_75t_R
XU218 n564 n152 N7 NAND2xp5_ASAP7_75t_R
XU219 n565 n149 N6 NAND2xp5_ASAP7_75t_R
XU220 cnt[0] n241 n240 OR2x2_ASAP7_75t_R
XU221 cnt[0] n561 INVx1_ASAP7_75t_R
XU222 cnt[2] n151 n150 NAND2xp5_ASAP7_75t_R
XU223 n243 N92 INVx1_ASAP7_75t_R
XU224 n245 N93 INVx1_ASAP7_75t_R
XU225 n247 N94 INVx1_ASAP7_75t_R
XU226 n248 N95 INVx1_ASAP7_75t_R
XU227 n244 n249 INVx1_ASAP7_75t_R
XU228 n246 n250 INVx1_ASAP7_75t_R
XU229 n251 N191 INVx1_ASAP7_75t_R
XU230 n253 N192 INVx1_ASAP7_75t_R
XU231 n255 N193 INVx1_ASAP7_75t_R
XU232 n256 N194 INVx1_ASAP7_75t_R
XU233 n252 n257 INVx1_ASAP7_75t_R
XU234 n254 n258 INVx1_ASAP7_75t_R
XU235 n259 N164 INVx1_ASAP7_75t_R
XU236 n261 N165 INVx1_ASAP7_75t_R
XU237 n263 N166 INVx1_ASAP7_75t_R
XU238 n265 N167 INVx1_ASAP7_75t_R
XU239 n266 N168 INVx1_ASAP7_75t_R
XU240 n260 n267 INVx1_ASAP7_75t_R
XU241 n262 n268 INVx1_ASAP7_75t_R
XU242 n264 n269 INVx1_ASAP7_75t_R
XU243 n270 N83 INVx1_ASAP7_75t_R
XU244 n272 N84 INVx1_ASAP7_75t_R
XU245 n274 N85 INVx1_ASAP7_75t_R
XU246 n275 N86 INVx1_ASAP7_75t_R
XU247 n271 n276 INVx1_ASAP7_75t_R
XU248 n273 n277 INVx1_ASAP7_75t_R
XU249 n278 N101 INVx1_ASAP7_75t_R
XU250 n280 N102 INVx1_ASAP7_75t_R
XU251 n282 N103 INVx1_ASAP7_75t_R
XU252 n283 N104 INVx1_ASAP7_75t_R
XU253 n279 n284 INVx1_ASAP7_75t_R
XU254 n281 n285 INVx1_ASAP7_75t_R
XU255 n286 N227 INVx1_ASAP7_75t_R
XU256 n288 N228 INVx1_ASAP7_75t_R
XU257 n290 N229 INVx1_ASAP7_75t_R
XU258 n292 N230 INVx1_ASAP7_75t_R
XU259 n293 N231 INVx1_ASAP7_75t_R
XU260 n287 n294 INVx1_ASAP7_75t_R
XU261 n289 n295 INVx1_ASAP7_75t_R
XU262 n291 n296 INVx1_ASAP7_75t_R
XU263 n297 add_1_root_add_0_root_add_96_31_A_1_ INVx1_ASAP7_75t_R
XU264 n299 add_1_root_add_0_root_add_96_31_A_2_ INVx1_ASAP7_75t_R
XU265 n301 add_1_root_add_0_root_add_96_31_A_3_ INVx1_ASAP7_75t_R
XU266 n303 add_1_root_add_0_root_add_96_31_A_4_ INVx1_ASAP7_75t_R
XU267 n305 add_1_root_add_0_root_add_96_31_A_5_ INVx1_ASAP7_75t_R
XU268 n306 add_1_root_add_0_root_add_96_31_A_6_ INVx1_ASAP7_75t_R
XU269 n298 n307 INVx1_ASAP7_75t_R
XU270 n300 n308 INVx1_ASAP7_75t_R
XU271 n302 n309 INVx1_ASAP7_75t_R
XU272 n304 n310 INVx1_ASAP7_75t_R
XU273 n311 N245 INVx1_ASAP7_75t_R
XU274 n313 N246 INVx1_ASAP7_75t_R
XU275 n315 N247 INVx1_ASAP7_75t_R
XU276 n316 N248 INVx1_ASAP7_75t_R
XU277 n312 n317 INVx1_ASAP7_75t_R
XU278 n314 n318 INVx1_ASAP7_75t_R
XU279 n319 N263 INVx1_ASAP7_75t_R
XU280 n321 N264 INVx1_ASAP7_75t_R
XU281 n323 N265 INVx1_ASAP7_75t_R
XU282 n324 N266 INVx1_ASAP7_75t_R
XU283 n320 n325 INVx1_ASAP7_75t_R
XU284 n322 n326 INVx1_ASAP7_75t_R
XU285 n327 N173 INVx1_ASAP7_75t_R
XU286 n329 N174 INVx1_ASAP7_75t_R
XU287 n331 N175 INVx1_ASAP7_75t_R
XU288 n333 N176 INVx1_ASAP7_75t_R
XU289 n334 N177 INVx1_ASAP7_75t_R
XU290 n328 n335 INVx1_ASAP7_75t_R
XU291 n330 n336 INVx1_ASAP7_75t_R
XU292 n332 n337 INVx1_ASAP7_75t_R
XU293 n338 N137 INVx1_ASAP7_75t_R
XU294 n340 N138 INVx1_ASAP7_75t_R
XU295 n342 N139 INVx1_ASAP7_75t_R
XU296 n343 N140 INVx1_ASAP7_75t_R
XU297 n339 n344 INVx1_ASAP7_75t_R
XU298 n341 n345 INVx1_ASAP7_75t_R
XU299 n346 N74 INVx1_ASAP7_75t_R
XU300 n348 N75 INVx1_ASAP7_75t_R
XU301 n350 N76 INVx1_ASAP7_75t_R
XU302 n351 N77 INVx1_ASAP7_75t_R
XU303 n347 n352 INVx1_ASAP7_75t_R
XU304 n349 n353 INVx1_ASAP7_75t_R
XU305 n354 add_5_root_add_0_root_add_96_31_B_1_ INVx1_ASAP7_75t_R
XU306 n356 add_5_root_add_0_root_add_96_31_B_2_ INVx1_ASAP7_75t_R
XU307 n358 add_5_root_add_0_root_add_96_31_B_3_ INVx1_ASAP7_75t_R
XU308 n360 add_5_root_add_0_root_add_96_31_B_4_ INVx1_ASAP7_75t_R
XU309 n361 add_5_root_add_0_root_add_96_31_B_5_ INVx1_ASAP7_75t_R
XU310 n355 n362 INVx1_ASAP7_75t_R
XU311 n357 n363 INVx1_ASAP7_75t_R
XU312 n359 n364 INVx1_ASAP7_75t_R
XU313 n365 add_1_root_add_0_root_add_96_31_B_1_ INVx1_ASAP7_75t_R
XU314 n367 add_1_root_add_0_root_add_96_31_B_2_ INVx1_ASAP7_75t_R
XU315 n369 add_1_root_add_0_root_add_96_31_B_3_ INVx1_ASAP7_75t_R
XU316 n371 add_1_root_add_0_root_add_96_31_B_4_ INVx1_ASAP7_75t_R
XU317 n373 add_1_root_add_0_root_add_96_31_B_5_ INVx1_ASAP7_75t_R
XU318 n374 add_1_root_add_0_root_add_96_31_B_6_ INVx1_ASAP7_75t_R
XU319 n366 n375 INVx1_ASAP7_75t_R
XU320 n368 n376 INVx1_ASAP7_75t_R
XU321 n370 n377 INVx1_ASAP7_75t_R
XU322 n372 n378 INVx1_ASAP7_75t_R
XU323 n379 N209 INVx1_ASAP7_75t_R
XU324 n381 N210 INVx1_ASAP7_75t_R
XU325 n383 N211 INVx1_ASAP7_75t_R
XU326 n384 N212 INVx1_ASAP7_75t_R
XU327 n380 n385 INVx1_ASAP7_75t_R
XU328 n382 n386 INVx1_ASAP7_75t_R
XU329 n387 N119 INVx1_ASAP7_75t_R
XU330 n389 N120 INVx1_ASAP7_75t_R
XU331 n391 N121 INVx1_ASAP7_75t_R
XU332 n392 N122 INVx1_ASAP7_75t_R
XU333 n388 n393 INVx1_ASAP7_75t_R
XU334 n390 n394 INVx1_ASAP7_75t_R
XU335 n395 add_6_root_add_0_root_add_96_31_B_1_ INVx1_ASAP7_75t_R
XU336 n397 add_6_root_add_0_root_add_96_31_B_2_ INVx1_ASAP7_75t_R
XU337 n399 add_6_root_add_0_root_add_96_31_B_3_ INVx1_ASAP7_75t_R
XU338 n401 add_6_root_add_0_root_add_96_31_B_4_ INVx1_ASAP7_75t_R
XU339 n402 add_6_root_add_0_root_add_96_31_B_5_ INVx1_ASAP7_75t_R
XU340 n396 n403 INVx1_ASAP7_75t_R
XU341 n398 n404 INVx1_ASAP7_75t_R
XU342 n400 n405 INVx1_ASAP7_75t_R
XU343 n406 N110 INVx1_ASAP7_75t_R
XU344 n408 N111 INVx1_ASAP7_75t_R
XU345 n410 N112 INVx1_ASAP7_75t_R
XU346 n411 N113 INVx1_ASAP7_75t_R
XU347 n407 n412 INVx1_ASAP7_75t_R
XU348 n409 n413 INVx1_ASAP7_75t_R
XU349 n414 N182 INVx1_ASAP7_75t_R
XU350 n416 N183 INVx1_ASAP7_75t_R
XU351 n418 N184 INVx1_ASAP7_75t_R
XU352 n419 N185 INVx1_ASAP7_75t_R
XU353 n415 n420 INVx1_ASAP7_75t_R
XU354 n417 n421 INVx1_ASAP7_75t_R
XU355 n422 N38 INVx1_ASAP7_75t_R
XU356 n424 N39 INVx1_ASAP7_75t_R
XU357 n426 N40 INVx1_ASAP7_75t_R
XU358 n428 N41 INVx1_ASAP7_75t_R
XU359 n429 N42 INVx1_ASAP7_75t_R
XU360 n423 n430 INVx1_ASAP7_75t_R
XU361 n425 n431 INVx1_ASAP7_75t_R
XU362 n427 n432 INVx1_ASAP7_75t_R
XU363 n433 N200 INVx1_ASAP7_75t_R
XU364 n435 N201 INVx1_ASAP7_75t_R
XU365 n437 N202 INVx1_ASAP7_75t_R
XU366 n438 N203 INVx1_ASAP7_75t_R
XU367 n434 n439 INVx1_ASAP7_75t_R
XU368 n436 n440 INVx1_ASAP7_75t_R
XU369 n441 N236 INVx1_ASAP7_75t_R
XU370 n443 N237 INVx1_ASAP7_75t_R
XU371 n445 N238 INVx1_ASAP7_75t_R
XU372 n446 N239 INVx1_ASAP7_75t_R
XU373 n442 n447 INVx1_ASAP7_75t_R
XU374 n444 n448 INVx1_ASAP7_75t_R
XU375 n449 N47 INVx1_ASAP7_75t_R
XU376 n451 N48 INVx1_ASAP7_75t_R
XU377 n453 N49 INVx1_ASAP7_75t_R
XU378 n455 N50 INVx1_ASAP7_75t_R
XU379 n456 N51 INVx1_ASAP7_75t_R
XU380 n450 n457 INVx1_ASAP7_75t_R
XU381 n452 n458 INVx1_ASAP7_75t_R
XU382 n454 n459 INVx1_ASAP7_75t_R
XU383 n460 N128 INVx1_ASAP7_75t_R
XU384 n462 N129 INVx1_ASAP7_75t_R
XU385 n464 N130 INVx1_ASAP7_75t_R
XU386 n465 N131 INVx1_ASAP7_75t_R
XU387 n461 n466 INVx1_ASAP7_75t_R
XU388 n463 n467 INVx1_ASAP7_75t_R
XU389 n468 N65 INVx1_ASAP7_75t_R
XU390 n470 N66 INVx1_ASAP7_75t_R
XU391 n472 N67 INVx1_ASAP7_75t_R
XU392 n473 N68 INVx1_ASAP7_75t_R
XU393 n469 n474 INVx1_ASAP7_75t_R
XU394 n471 n475 INVx1_ASAP7_75t_R
XU395 n476 N56 INVx1_ASAP7_75t_R
XU396 n478 N57 INVx1_ASAP7_75t_R
XU397 n480 N58 INVx1_ASAP7_75t_R
XU398 n482 N59 INVx1_ASAP7_75t_R
XU399 n483 N60 INVx1_ASAP7_75t_R
XU400 n477 n484 INVx1_ASAP7_75t_R
XU401 n479 n485 INVx1_ASAP7_75t_R
XU402 n481 n486 INVx1_ASAP7_75t_R
XU403 n487 N146 INVx1_ASAP7_75t_R
XU404 n489 N147 INVx1_ASAP7_75t_R
XU405 n491 N148 INVx1_ASAP7_75t_R
XU406 n493 N149 INVx1_ASAP7_75t_R
XU407 n495 N150 INVx1_ASAP7_75t_R
XU408 n496 N151 INVx1_ASAP7_75t_R
XU409 n488 n497 INVx1_ASAP7_75t_R
XU410 n490 n498 INVx1_ASAP7_75t_R
XU411 n492 n499 INVx1_ASAP7_75t_R
XU412 n494 n500 INVx1_ASAP7_75t_R
XU413 n501 N155 INVx1_ASAP7_75t_R
XU414 n503 N156 INVx1_ASAP7_75t_R
XU415 n505 N157 INVx1_ASAP7_75t_R
XU416 n507 N158 INVx1_ASAP7_75t_R
XU417 n509 N159 INVx1_ASAP7_75t_R
XU418 n510 N160 INVx1_ASAP7_75t_R
XU419 n502 n511 INVx1_ASAP7_75t_R
XU420 n504 n512 INVx1_ASAP7_75t_R
XU421 n506 n513 INVx1_ASAP7_75t_R
XU422 n508 n514 INVx1_ASAP7_75t_R
XU423 n515 N218 INVx1_ASAP7_75t_R
XU424 n517 N219 INVx1_ASAP7_75t_R
XU425 n519 N220 INVx1_ASAP7_75t_R
XU426 n521 N221 INVx1_ASAP7_75t_R
XU427 n523 N222 INVx1_ASAP7_75t_R
XU428 n525 N223 INVx1_ASAP7_75t_R
XU429 n526 N224 INVx1_ASAP7_75t_R
XU430 n516 n527 INVx1_ASAP7_75t_R
XU431 n518 n528 INVx1_ASAP7_75t_R
XU432 n520 n529 INVx1_ASAP7_75t_R
XU433 n522 n530 INVx1_ASAP7_75t_R
XU434 n524 n531 INVx1_ASAP7_75t_R
XU435 n532 N254 INVx1_ASAP7_75t_R
XU436 n534 N255 INVx1_ASAP7_75t_R
XU437 n536 N256 INVx1_ASAP7_75t_R
XU438 n538 N257 INVx1_ASAP7_75t_R
XU439 n540 N258 INVx1_ASAP7_75t_R
XU440 n542 N259 INVx1_ASAP7_75t_R
XU441 n543 N260 INVx1_ASAP7_75t_R
XU442 n533 n544 INVx1_ASAP7_75t_R
XU443 n535 n545 INVx1_ASAP7_75t_R
XU444 n537 n546 INVx1_ASAP7_75t_R
XU445 n539 n547 INVx1_ASAP7_75t_R
XU446 n541 n548 INVx1_ASAP7_75t_R
XU447 n588 n562 n598 NAND2xp5_ASAP7_75t_R
XU448 input_buffer[3] n561 n567 NAND2xp5_ASAP7_75t_R
XU449 input_buffer[4] cnt[0] n566 NAND2xp5_ASAP7_75t_R
XU450 n567 n566 n600 NAND2xp5_ASAP7_75t_R
XU451 n600 N6 n571 NAND2xp5_ASAP7_75t_R
XU452 input_buffer[5] n561 n569 NAND2xp5_ASAP7_75t_R
XU453 input_buffer[6] cnt[0] n568 NAND2xp5_ASAP7_75t_R
XU454 n569 n568 n621 NAND2xp5_ASAP7_75t_R
XU455 n621 n562 n570 NAND2xp5_ASAP7_75t_R
XU456 n571 n570 n612 NAND2xp5_ASAP7_75t_R
XU457 input_buffer[7] n561 n573 NAND2xp5_ASAP7_75t_R
XU458 input_buffer[8] cnt[0] n572 NAND2xp5_ASAP7_75t_R
XU459 n573 n572 n620 NAND2xp5_ASAP7_75t_R
XU460 input_buffer[4] n561 n578 NAND2xp5_ASAP7_75t_R
XU461 input_buffer[5] cnt[0] n577 NAND2xp5_ASAP7_75t_R
XU462 n578 n577 n607 NAND2xp5_ASAP7_75t_R
XU463 n607 N6 n582 NAND2xp5_ASAP7_75t_R
XU464 input_buffer[6] n561 n580 NAND2xp5_ASAP7_75t_R
XU465 input_buffer[7] cnt[0] n579 NAND2xp5_ASAP7_75t_R
XU466 n580 n579 n630 NAND2xp5_ASAP7_75t_R
XU467 n630 n562 n581 NAND2xp5_ASAP7_75t_R
XU468 n582 n581 n616 NAND2xp5_ASAP7_75t_R
XU469 input_buffer[8] n561 n629 NAND2xp5_ASAP7_75t_R
XU470 input_buffer[0] n561 n587 NAND2xp5_ASAP7_75t_R
XU471 input_buffer[1] cnt[0] n586 NAND2xp5_ASAP7_75t_R
XU472 n587 n586 n593 NAND2xp5_ASAP7_75t_R
XU473 n593 n562 n605 NAND2xp5_ASAP7_75t_R
XU474 n588 N6 n592 NAND2xp5_ASAP7_75t_R
XU475 input_buffer[1] n561 n590 NAND2xp5_ASAP7_75t_R
XU476 input_buffer[2] cnt[0] n589 NAND2xp5_ASAP7_75t_R
XU477 n590 n589 n599 NAND2xp5_ASAP7_75t_R
XU478 n599 n562 n591 NAND2xp5_ASAP7_75t_R
XU479 n592 n591 n613 NAND2xp5_ASAP7_75t_R
XU480 n593 N6 n597 NAND2xp5_ASAP7_75t_R
XU481 input_buffer[2] n561 n595 NAND2xp5_ASAP7_75t_R
XU482 input_buffer[3] cnt[0] n594 NAND2xp5_ASAP7_75t_R
XU483 n595 n594 n606 NAND2xp5_ASAP7_75t_R
XU484 n606 n562 n596 NAND2xp5_ASAP7_75t_R
XU485 n597 n596 n617 NAND2xp5_ASAP7_75t_R
XU486 n599 N6 n602 NAND2xp5_ASAP7_75t_R
XU487 n600 n562 n601 NAND2xp5_ASAP7_75t_R
XU488 n602 n601 n625 NAND2xp5_ASAP7_75t_R
XU489 n606 N6 n609 NAND2xp5_ASAP7_75t_R
XU490 n607 n562 n608 NAND2xp5_ASAP7_75t_R
XU491 n609 n608 n628 NAND2xp5_ASAP7_75t_R
XU492 N279 n549 INVx1_ASAP7_75t_R
XU493 N278 n550 INVx1_ASAP7_75t_R
XU494 N277 n551 INVx1_ASAP7_75t_R
XU495 N276 n552 INVx1_ASAP7_75t_R
XU496 N275 n553 INVx1_ASAP7_75t_R
XU497 N274 n554 INVx1_ASAP7_75t_R
XU498 N273 n555 INVx1_ASAP7_75t_R
XU499 N272 n556 INVx1_ASAP7_75t_R
XU500 N271 n557 INVx1_ASAP7_75t_R
XU501 rst_n n558 INVx1_ASAP7_75t_R
XU502 n617 n559 INVx1_ASAP7_75t_R
XU503 n613 n560 INVx1_ASAP7_75t_R
XU504 n242 n563 INVx1_ASAP7_75t_R
XU505 n241 n564 INVx1_ASAP7_75t_R
XU506 n151 n565 INVx1_ASAP7_75t_R
XU507 input_buffer[0] cnt[0] n588 AND2x2_ASAP7_75t_R
XU508 n620 N6 n574 AND2x2_ASAP7_75t_R
XU509 n598 n242 n604 AND2x2_ASAP7_75t_R
XU510 n605 n242 n611 AND2x2_ASAP7_75t_R
XU511 n562 n629 n632 AND2x2_ASAP7_75t_R
.ENDS


.SUBCKT CIM_adder_tree_DW01_add_1 A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] CO
XU1_7 A[7] B[7] n3 n9 n10 FAx1_ASAP7_75t_R
XU1_6 A[6] B[6] n4 n11 n12 FAx1_ASAP7_75t_R
XU1_5 A[5] B[5] n5 n13 n14 FAx1_ASAP7_75t_R
XU1_4 A[4] B[4] n6 n15 n16 FAx1_ASAP7_75t_R
XU1_3 A[3] B[3] n7 n17 n18 FAx1_ASAP7_75t_R
XU1_2 A[2] B[2] n8 n19 n20 FAx1_ASAP7_75t_R
XU1_1 A[1] B[1] n1 n21 n22 FAx1_ASAP7_75t_R
XU1 A[0] B[0] n1 AND2x2_ASAP7_75t_R
XU2 B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU3 n11 n3 INVx1_ASAP7_75t_R
XU4 n13 n4 INVx1_ASAP7_75t_R
XU5 n15 n5 INVx1_ASAP7_75t_R
XU6 n17 n6 INVx1_ASAP7_75t_R
XU7 n19 n7 INVx1_ASAP7_75t_R
XU8 n21 n8 INVx1_ASAP7_75t_R
XU9 n9 SUM[8] INVx1_ASAP7_75t_R
XU10 n10 SUM[7] INVx1_ASAP7_75t_R
XU11 n12 SUM[6] INVx1_ASAP7_75t_R
XU12 n14 SUM[5] INVx1_ASAP7_75t_R
XU13 n16 SUM[4] INVx1_ASAP7_75t_R
XU14 n18 SUM[3] INVx1_ASAP7_75t_R
XU15 n20 SUM[2] INVx1_ASAP7_75t_R
XU16 n22 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT CIM_adder_tree_DW01_add_0 A[12] A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[12] B[11] B[10] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[12] SUM[11] SUM[10] SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0] CO
XU1_11 A[11] B[11] n5 n15 n16 FAx1_ASAP7_75t_R
XU1_10 A[10] B[10] n6 n17 n18 FAx1_ASAP7_75t_R
XU1_9 A[9] B[9] n7 n19 n20 FAx1_ASAP7_75t_R
XU1_8 A[8] B[8] n8 n21 n22 FAx1_ASAP7_75t_R
XU1_7 A[7] B[7] n9 n23 n24 FAx1_ASAP7_75t_R
XU1_6 A[6] B[6] n10 n25 n26 FAx1_ASAP7_75t_R
XU1_5 A[5] B[5] n11 n27 n28 FAx1_ASAP7_75t_R
XU1_4 A[4] B[4] n12 n29 n30 FAx1_ASAP7_75t_R
XU1_3 A[3] B[3] n13 n31 n32 FAx1_ASAP7_75t_R
XU1_2 A[2] B[2] n14 n33 n34 FAx1_ASAP7_75t_R
XU1_1 A[1] B[1] n1 n35 n36 FAx1_ASAP7_75t_R
XU1 A[0] B[0] n1 AND2x2_ASAP7_75t_R
XU2 A[12] n4 SUM[12] XOR2xp5_ASAP7_75t_R
XU3 B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU4 n15 n4 INVx1_ASAP7_75t_R
XU5 n17 n5 INVx1_ASAP7_75t_R
XU6 n19 n6 INVx1_ASAP7_75t_R
XU7 n21 n7 INVx1_ASAP7_75t_R
XU8 n23 n8 INVx1_ASAP7_75t_R
XU9 n25 n9 INVx1_ASAP7_75t_R
XU10 n27 n10 INVx1_ASAP7_75t_R
XU11 n29 n11 INVx1_ASAP7_75t_R
XU12 n31 n12 INVx1_ASAP7_75t_R
XU13 n33 n13 INVx1_ASAP7_75t_R
XU14 n35 n14 INVx1_ASAP7_75t_R
XU15 n20 SUM[9] INVx1_ASAP7_75t_R
XU16 n22 SUM[8] INVx1_ASAP7_75t_R
XU17 n24 SUM[7] INVx1_ASAP7_75t_R
XU18 n26 SUM[6] INVx1_ASAP7_75t_R
XU19 n28 SUM[5] INVx1_ASAP7_75t_R
XU20 n30 SUM[4] INVx1_ASAP7_75t_R
XU21 n32 SUM[3] INVx1_ASAP7_75t_R
XU22 n34 SUM[2] INVx1_ASAP7_75t_R
XU23 n36 SUM[1] INVx1_ASAP7_75t_R
XU24 n16 SUM[11] INVx1_ASAP7_75t_R
XU25 n18 SUM[10] INVx1_ASAP7_75t_R
.ENDS


